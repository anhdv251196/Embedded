XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��.���o4VB�F$\��y�s����H�V	$�ȫ����q K4�a�H;>�0?�[�*�ۓ�����Fe�P����I�rΩ�9���2h+�E�xl�p�mUot����H~`��F�^��}�Y5�f�
(�٪I��o�m,�q��c�]ϙ�"���Ǻ1Ln�)OS�xm��:���� �ݖ��9c���ĭ4���9g+�6_�Ĵ�����t���B��6HO�ߜg"q:<$
1o-Ac�Y�`��<-�x܋r^��K01�5J�C�>���;�b���f ]W����c�[�a�5�hǪ��u6��
p��2�f�� �n�ea����Ka�}g�.6���*x���s~����N���R�����H)~Z�x�?�ӱ�J��9�/+0P
�"���}�}wgIW���̋�����up:3�Xl� �dpć�P4
�-L��#
�ʣ��:H^�X	i�0��-� ���a_�|XW�HS-�/湼5��AK+[x��-J#�t)��W��=�-�k�vWY!*�B��'��V1Rz�W	ռ�y�34����}͙"I�ӎ�VP�x��������-�m��9�ڦ�qwBÆ��z�+�Ճz��U㫪V�ռm�ZH>ʨGM�SR�n����N��i����Ca�
K��[�}�Uٻ�*BSS+����g�EȀlR�k8Q�i	V�!�bɐB�!w��!��#2��,�4�a��L���M�.�a=��8�iu'Q��Ս���jy���=�~��� � XlxVHYEB    1ee7     570[�#dΖI�q��wpW��FV��v�W�����<̔��'9�zk+T�kS�MN��L�a�Q�4��b��(�c��/s{[��$g�v�Fw-U��ο�:�'�p[_y!�,fO��,�J������A=H NG�3݄Sk�]���м�"�	�'�t�~y�"@��-4g F���_H���
����_��g�<z}����NoNv�RBCj��'^a�c���v7�#۫]��o0��v�L�@�_${�؏A#ɺ�{f���'ګ^�Jz�o�	��A�bpk �t�=v�.֒�Hv��!��14O���^��?u�`�U3\�P��@ގ��N&^G�MK��1hpy��`�n��a�������J�C�(���J�sS�q�v��!z ��/~<⁝�unj�)#���b����t�(V�#��"9�f�֗�s��R����!�����U ���\ �'���E��l�[��mE�i����F�@����\Z?.��z��Z��M���S�_�kԣ�%�oK��!��ty�b���� 3?���]l�	a8}S��Lti41��J�� Z��y{�����R�E�:�zY��شc�q�8�[4!�|�GK��P�$6�й>?��/8��Q�aX�f<	���7�čs��ν��6[#�,]���f�{$C9��C>�hj\rG����E��.ʺ�5@�y�ЀDI�y��/�3�zd��k�F;aN��'���н9 2ßנ���V�0����C�Y�E�C`Lq``n����R��#�������e�<��Rt>^u�*#�
��u*"�A��زU]�/;;$��<w�2�x��n��I��3i��g�2=�F�1N����|���<�=7F��׈�6{�¸�e������Aۑ�ϵ�U�~^F�q�Cf��G��g	�VD���jZ;v�Ec��؉��x:�}�5-X� ����'�_#�v{�	W��v�:�~�u#q >�}v,Z��,l�]F82�ḃ^�MV�y$h���_�s�NM[�u�k��AEa��Ő�� !Tz�2��a2�ዕ�e�;�������Cc�M�0%t���Ms��ϋ��DReGӮ��&��]Q�h~@$y,K��=�xz茏N�[$�$�����l�T���£����+NѪOd�j���:>���x� ���£����h�_s�U�:�g��T{a��ظ���� wz�1.L`��3H��Ү�^1�[�o ڎ$<��c���~)���-�eJϥS��-�Px��Dq�pj_W�t�֒}��F�[L�Cݶ�I�x���ɕ�3:�e-ѻ�����+�m7��<��k��=�$���ϓ�lg3��5.h9�E;EK��d|��