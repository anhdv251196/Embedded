XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��LBn��Eu>ʯ��ti�\��:t�r���TK�®���V��4�����P�׽��zcȪ�ʿۺ�հ�um�q�݂�-_#�~�ɒ��>2C�G;��I��z�������k���_�_%�<���2��O���͸�M6���K�����n
!�F"?�0v�zxߡ:�|���4
�s���4�	R609��:r��!^�,W�5$r��1@\$�*���?��2k
T,P����%�3�X�b3A����K��b��ןG�g��4��.�	�xa�L�4pSrE�L�x�}��?H�L�M(81�� S<�󌷑���dc��+�./k�фW��G�V3�O�t��nٍ�bN���
�aQH�������@@� ���g&�;�F��T95|���:J\����0U)H�%⟂�由���xkP/�e`w_�I��q�CW��C#�H*詹1y8�$�j����H\K�D~'Uդ��\��F�&#�F^�r*��w�I�c�%Q������(�;	��nOw�������fƲ֘���O��dϲs�n���ښ����g���fbY�^��6�I�l����ם
Ė=\���.�ARi��Ua������0ZL���M_*�(��t\���Ł�]��S9�Ө\��F�V?q�.���m@��U�@���w��������q��L��R�����(��W�y��a�;/�/���bߥE�|~��k/���W>����s;����XlxVHYEB    5ff4    1040����N/1���KՐ�,��ow�&���)"�p�\fˍ5E_�!�	)Ct�g��������Z8�['��\�tQ|}"����q-�`��>}xbٸ����6_I�V���:iT��m�@��X���3ik2�_��,D��FP�S��xz��r�ܵe�I?͘�ú��)2r\^��✔i��9%<D��o�q�fc��-�\ټ�=3>����yU�Fy@o|N[��LyGK��� ���%����#y��h���{]ѹV��(��b�MA����^���#�n�R��-bU�)Rz!��(�p]<��нmP���{�<��"��nF��|�T���ؙI�z[CT��Vޱ����LY�ę��h֐j`܉¨��)�Vs����3'��eԄ��^�/���g����'E&���������%����ڠV�yƨTG������s�^5�7��nQP��r�!�L��x͒������Ȍ
�ӄ�CW���C�<x-pċ��ﾪ�sw�B����V׺R�RnCK(�%�,sl�}�%$�>���jݬ����O��7e�k@9M!����
�A�#B��i�aLp�ldEYU�Q����dR`ܦxQ �����{����{��(E�U�#��j4r:�Q�طa<��j�FD+���&�Q7��K�R�(C^���Zk~;�N�P��k�.�EgH���� ���k.�HPc�'�Dzj�ߢ�Cgi�p�SV���wP.��t�*��jv�[x���,o�0G���F��C���������c��A�%�>�I�+�s��J|�E(R�P"�30 ���J����5��7%�"�N�Z�[)������Mr=�Z��6�t6}�A������_/�3���̹0Ϫ5��zZ��@������9��p5a�"	�u0䌶`�����=��ث(��DȌ �~�:��]�m��֢�Nwa��΁��-ɔ��[u��d�g&�����%?<�6wI��Ő��z�˫�� iw1��I��mj?=��r?^��u9(�4[tJ�ȟْ����YF'����X�Z��	t^%��O���0�q���m{d�T�Eyɚ{�x��͘u��@t����c{���c�T~9r���fyY�����0���\�S!�'k^�ʨ�k�j]�_�½� ��B^4��˩p�(��ݞF��} lK�1%���EU��.%Jb{��H��Z�F��W��$gn�A���k0-�7� �=?�
)���W��
���+�Z���6<X���l~��5g9�+ɢp	54��sU�[���O9��:v��������w��}������O�M"��vW��#��Jɸt�� �Wu6�7�%C�0�Z�m����_k{/),D�����n E8�ִ\ڷo����SN�;�Q�|��!GK�	 ����A��A��7[�ܠcL���~T(C@1mF�֦�;��5X�$�ce���:�j<߳�i���k�r%J�q�yÿ�ߌP��[\�%�G�A<3�V9�_�Z�T�����/w;x4���4ʞg�������?�a��Gh+�+�W�������$[�qoy�l�c=ne)'���u"��i��7*YrȎ
P��{B�->��?�Əz��h���5KE�q�j�����ߺ'ب�#�eC�\C�SA�O�cwȦ��A/���_�ר�-A���<��
��b��G;ѕW�ɢ=V�뒤6�� #�@�@�ꯧ���|@�����=�\����^��j&���5�)��� �Z~.*�<�r�~0�6Q�U�褸�ğ�����f�Y�)Zo>�&����~����,��w�c��UZ�ے��u������^������Ad�]�Q�ykUsD ��r��������.�6�=�@H+�ƞɦ���h8�^��EHT9+��$�ѓ$_n�f)v-�M�\��
s<�}du��|h-���n8��Їʤ<�؀�͋#���!q�}_��.ЌH����NS��i܈������	�n�����^#�5I>���ܧ�҄��f��op�ZFh��^��89��ʰ�,����U�"�<����̨$����n?z����S��fds��=� Z�B�7uO�U�ry�˩ĶӞ\���L��h8UT9f�|�-�HL��ORX:{�U�i%S��r� <	�%��rH$��ᨘ��H;�l��Ս�Yr�:��	�6��}��i61{
Z�rl#CK�c��Ƙ�n�s���)Ӓ=��ޯ
��`�Hb)k���h�
H�w��a�B������<�Ā�����
�"���Px~�8
j&!ʿO�p|���'��fw�ɼ���qpq�T��VO�v���:�&��,����(� l�v���W����?`P�g駚�r��s�	= g  ��;ߑ��Ԍ#9��f�-��  �gݖ
^�܃�+k^�0=E!t�}��Qp&la��v���_`��Z�����B�0�xԮ�/ Mt�?{G�����Y��j8b�͎ܤ�U��'�F1�A��	l�� )�B�33 EUVd�+j����v���V#���Yf�����P�ʩ�⃟5s��n������=�R�͋��rJV��A/gԚ=8OI���0e�u�pR��(NQE��q��cȢY�P����YEG�Jx� �	G���L���e�ѽ���}���(d�E��?L3r��g)C�s]Q�e9��x��Y;l�g�C��C_)ê�Yx���tPme:�qL�n�
�T���ĥ��f��\FХ�*_���&�?�t�8��\L,+��G#~TZY�[�N�,{�7�Ju>n?	� (�D9s ��|��:���֯k8�E�Qg`�죹5�B3���W�P��@�����O����}��m[A�c�~�. ����@aB���7H��������ss�v�vЫٮ�/]�A�0� ���S֓WDz' ��:8,>��ԥ�s���
R�w�
�A�����[1AJE;��u��+O��"U�d�^+Ջ�S&!�W\�O&�N�8S�k����H��M VZ�,�~Q
?y�돰ᬑ$[��<�:g���zf[bכ1HG� M�S_	%����B��E��ԩD����c;�h��°�
���E�M[�p���ϊ=Sw`{�!{��։L`�`6�,piAA��q�h��6F;o����S����>B4Hh]��v�'b�}����N��:��`C9���㚺z�}�ȼ�o�W����G^"�I`Y�uSɫ'� �RJ��pI�꛲�$�v�V�1���PTr���|S�RJQ�u�V_�@�.j�\3�I��+j���u;�K���X�u���V���C�֋?�ˈ�n "f�+�^�:8l���n����8|�x�޶�u��$����+���=���C������b^���A3��l!�V�	��të��a>���6��j?�2�9��5�Y�k���hǤN��#��-���H��k�`+�{g�1|��r@t���J�=��L��B��]����
�g2��%TU^ŮC�����ޤ�ɨ�`�4#h�ou�k�E��^?�q�����M��.o�Y{3b�p9���NÂ�GL�R�+��Cp�-=�9�Z��0��mN���"�������wƄ�����.��!�F!�D�eX'���.���>���k
�7�f�f�^A��
����X+hN n�P)�~���y4�Qd��� ������@Y���F��o���Ɍ���?�>>_��j�A�>(��7�9�f�';w�g�����ڙ<�� e	���@�q�$�&)��=��`�/�3��*���Z����`�g�1M��m/]r[��B�Va�둇����s0���(�>@2�,Mۑ��S�2-�[в��=�I{
��Z���.����5�Hn}�y���u]��g������������4Nk���`�v��ܧ�%s�TЀ��sz&�N�tB�)� VeW0}�^�����b=�
���
��d�0��&��~ըu�϶���zfZ�#����'��;�9=Ǐ9�ӛYy�H*�i�F��6^���z*�d)Ԃ}&7��	q�R����K\h 'A��L�ݾ�*Sjm�l��Y߅�F�ӡ�wۀ��DN/�UN���/|O~�Sz-BE�+3$