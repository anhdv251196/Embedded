XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��;�DA��Z� ��A�S^N��/��Բ_�Y��Px�������X:)*�V8������FFМ�?21�Q��*����]R���]��hʣ�6��)�r�����y���n��coU�z=7p�V'��d�h�Vx�T1���_L��h1���|@Ҫk_�H�n)ڐ�sgi�݌�qs!�1��k���-��B�#.�����Y������(5�S���h��R���IU\��I\8�w[޸	�����8�f$<�����C��*m�4R�
����Z�o]���ď yc�����"+��t�������_\�z�1X^�/���,W;r�x贁�5_�8@�k']�3�m�V�d�b��<h�2�����eύ3:���,���}b&��O�L��j���QS��7u��h���
g�I�Gi�O��w@j��&� Ξ>
�t��5�D�KuAS3(��m	���,9t�@�����i;�
K�� e�����{��=XP���-�⟈{)�3B{��S���/d��9�
*�Ui+VsO�u*����zw��z�8��G�)�{'���(�|x����a�ot�3#F$\�b��ƻ�<x�Z�L�Ut�o�٥�N�%�^��T_S�%����3#��P0�t'Nn�26=\9����+2���rVg�@'�#��T��?�e��r���c�>���_?�.H�Cw,����UOj��&��Kʯ�p���S���d�U�k�~��D�j��_� �2��q'P�e��{WP�=����D�~�XlxVHYEB    1cf8     790T���#X���w�Y{r��b�ر-�8�a�c�8��|�㇅��\���P0��ڴWOR����A�{����-���2��S>	s�����q������V��]����UR?�����"�)AF�ϊ�v4+J|�ղ�犏U�TL[��ާ�A�SIՀ2��,J��	�!q+�r��s7Z�[�����:�>���R�����m�5I�NӼ��N�0�VdUa�F<�)i\��f`A/��]`��p(�%�gF�F��qUkf�W�|񣶈��Ϯ.�|��X�*q���}|�2}7�w�'��AB%k$��m��X���	$�j=�p��o�E��8 E&�ߧ��[�g��&�{\���?�p�����D��#'������K
)�ean5�.~�l��	c�f��>;����Ou����S���/W�!`(��ëK\}�<�J<���̮�%�5�����2�I����9	x�lnk0���+��-���!�����s��c�&�qS3�Z�rm,ta��%�ŗ_E�ч{��w7��^L+�7kH)3Z�R����e�z�Z��M���A+��4RZ�$�L	[�������$ԩ�T���<�,chñѸ�r)`@"��_٨#Aݚ-���4��Nz`���.=��Y�\X�1�����?},�I�_�*[�J�A[~���E,t���d����a2����^�wX�5���{#�)�(�3K���&-�^��_C�0\vt�q�P�>$��ٚ0�>��餹#�ޕn:o�+y֫��P�n��v#5�l#�#v}e��ʠ/�I�S�B.db�сĕG� h�kS����Y�1$�%p����ԗ�zU�A��V��w�[wo݂�gJ��营��i�0�����a�v'�9^C��btK� �j8���hFO%��̟Q�����N�P��h�VܹEta���f>��m�ʼoq= *� ]�%��'��ѳp���Ÿ�X��0_�l)�k�l�eu�&])��KY�J����ƴI�1�̸�;2�����pQv��j��8��O��f��`����J~y0�k�jV�v��l���5�u�?@;d�Ȼ|j��,�~5���9�v_���Q�H�K�s�y��.� Ɣm�?l~��a I��6��{��_��6�@��?��=�!Q�Zz��1/����B^���(d~��~��@6&�Q����`��
��3��_3���ը'!����+o���W<��A�@L�)8�G��4�9\���H*|����oLK���p���7�Ͷ���`�م���T������¾AU��/�?(Z�����껷s��P[B�9�0�$�Zy�7�U�� ĵt}y�0�p"֥�Y��5�J�Yr�=(�Է�i�r�AG�bc�Y3'��7�K�տd"�WZ����b�C��<��v��,ɒ��J���YC�4�1quHI�}˅���YL�8��w��!b�>7���[(���f[�ĝ�GP��x���K�!,���kl)@��	G�^�f���/�jm\ލ{1L/�+lJݢ�`a]e�+lx��J�5�m��g���@� l"�<�C��[-��q�I���(��A��(p��������% �uWl�Iv�͡�����Ԥ� 6x��
�ѩZ�LŚݡ����[y�Y�&�����	�QFYW��&f�;v���}?�pl�*�]�X�H;�C��j�O��Z��B钛y-��L��NLf�$�c_���,�:�hՃ�(B��a��.�Ѹ���kl�R����+�C�R:�og{��	�$oiP#�I��׆O"��'Z���>�&%d#��𗲵B�����{r�\�T���=%���齪�6�Go��f��Ɋʘ�l���+j��Nc���UA��|h�	�ڮ�5�r[���F��Ą�GXk�E�E�٠B���M�9n7w