XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����+�J��x|H:aXk@�<�(��qٲq��Vst?�Aeҕ��6{�1���:܇|�RѲӤ�_���@���ض<�v�f�h�j���^�	��Sw�C���	��]�����<.�;-x&YdEr�]1�w���5Xu��a	�PMM]�K-b31�fH�s�ג� �j����z�l+s0�϶�n(t�~9H5p��I�sr�~g��m�g�q=I`I��2L~�⍞U+CJ�������U�>���Y��  L!w�x�]j��okf����5F:�����)���P��oC��k�����TA�q-����X���b[�L�\j��]�j7�]�5K�8���Pq
��>z�1y������8�'D-���]�BV*Xі�'���M�֍F����@��vF�O��x4" Rdh0�5o�T�.�:_f�<)ZvR�ϯ������x3�D�?����@XR_r$/(|w�WSw��vBG�|َܸ+�N+�a���G�.(��d�dh�,u3����魂۝0��/2�k����3[�kI|z_�~PG��P[��'¼�DU_+�xK��=����:��-��o��+�4<������~sG�% V���3j!ϗ���E�O+�~�����uc>L��$[��E���q��6��V4�^͎� 4�N/͚,�q�O��l-�{&�s~�]t̒Ǣ�rea�Ec�،b���K����u��Y�LTO-�	�C!������᭕PȬp���XlxVHYEB    1578     5a0�̷����1��!9ew3�B���f��?�:6�69�50wwz�q)�	�ljy���'_������W�����5`�-�ݶ`e��.�w}��LA�jh�z^����F����}rp���-UW�s�0{���p:6^2��Z��#ͮbV���z��J���C�]���v	$�2p"Hw�s�#b�[�ͷ;����Y�U؆�`'���?��fWv�B����\ڑ3ăgy7j��0�j�8T\@�1)V��q�ah�u������U׊�&��io��a�1)�J ǈ�$G�e�M���ӵƺ�8�D̤(�A~)Z����\�2b�]'A�Ŀ<�L��{1KJz!�`8�����}���<H����b��)noT��S��ޓ��Sz,p'ЬuKW�0���R�}w�L�u��/@%��@�)�ō?��tx��:�}z��VuI��Ň�$ZB��9�d�#��%$���_�f}"�U�,4���f^K1��~ܸ�&��$�@���$���ө�Q�������-�{uhIc�0�
�+Ӄ�����S��F5f3}⟇�;i�H�t*�A�Ci�}T�6�d�y3��4hn�B5����5lyQ���-��c�e����˷�����0x$�#8 �L4�/�F��,�`�����;=��1�IZ�a +�$�<,QZ�qj\���dփ׬"v�\���V[\cf�-f3��ٜc^w0 ����
��B�^��R]#=��F�~�˪�6�J�95c�Z���'X}�'S!��7�ԀD�֪���*��D��xhu��xcA�[i��z�����K���	�u7��:^/��ڐ�Y���f�P����8G�H�`���&��#�I^n*ߣ���BQ�0�L���Ǹb¶���[%?�)��F��D��2&~��gI��SE�8G�\A�����J{�����J�l�Q�&���g�+���]��?�k(���Y�k2��dM��]�/~��:�)0��8#?/��7��:�������~��ed 6��吞V��U�Ww�v�vT�ܞA��X�-����3V("4O����t�B�N���|�c���.���Y�m�T_�9�����ʢ?DPK�f�Z�ͯ��z|��{I�L�k�=
7���ӰNߢ5�eR�Y�>+8�0jYX�DY7��l������f9�5hO9����J�226	��"��n�So�/n<w��Q$&���n�T�ٓ)VX�/2L'U�f��ƣL	�������YN/�<K2�J��y>�<oP;��R��� *�G �+���$��r0 �@�J�X�p$?�i4-JAf-���IZ9XI/��L��d�r���%��a�V�t�{2'�Gv$#X.�о8�OA���G��t�bb��0V���/?t����_X�f����Gj�0��;�����>��px\