XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��0���9f��~y?����ny<`�S�M.��.�=tc���m�C��OnŖ�\&6h�X�0z��EȞx��=B"��ݓ/���h�[9�;�5��\���'=,oX�2ʹ5�g\NpqQ�%�|�y�vE>z��H���GQ ��dw�;B�a����V����p�Wz���[��-e�l�4-��Tb-[&IV+i7�qS�dkr}��r]<�!�?'x���� Ŭa,�O�t��f���'���b��]t�N�X�0�<z-�2�Jd/��2���w��NhQ��i�e�QO��E$Ul\���c�YY}�k���lr@�3��Y�$��7j[G�N3��A��M��7T�N d�Y��8�~���/Iv1��9$f����0��y�������_2*7�wmlҢ�wC{�*�~j6a{� �§qn��܁����2�@2�֣�Z�����ÓQ�D��`�a��'H�y���p(Q����8"����Lǵ!��Z�+�5���8>&6 ]-���n���1>������U&�nv�s�c�gp���#b�\D�^��OUf̒L�4�B��ϩ$��FD�_;(�3�	��K�`���W�_��R���W�����:�!'�'�}�b?~��Y�n�Q1�����R���qW�)�25��6�*&-e�;y���n�(������Q֍�xpyrQ���5&~-�KR�Qk| ���J�|���)6��S'�F���I
�V��*V�E������w�<�WYM�b?n�|Ě��	�wH�5�XlxVHYEB     b88     3c0K(i�ʝ�6E"v?v�
g�
c�6.ql���5�9Q딦���et�"������k��j����J�,P+D���`��9�Zc\�	]^�N�c���DĒ���8'\��~�`��Q��_C_t��ds���tC��J��8�B�8��Ӗ��w���ZIm�a�ט�)t�����IՌ��%�u?�`�22�`�c��ղ��9�~���*FQ=A����5�_��*����v�%������{2�Ա�ѰH$G��&cx3�W^ � 5��V0�=�VC6ϰ�y��P���f3OS�b�h���mj^�//s%�����j�sD��bm.��Gg��$����"��|�iC���Yv�:hD����&���=�2�)��=��0ԕV3�˜��0bI�����w�%��S��ܿs�L�n���)�t�2�{�i���l�=]Ga���Jk�����EF��bF.վ��L�04��@6��9�R��z�)C$|8C&�(ț��$
����Jl�9�����A�݀��/�����X���P+���f�3��r(�)�Gx��K��gt���E�1C��M�F��$@�Y0Xm
���W������["�!�����\�8�$�;?H �Qm�L�=�\��]u���'0��O��9� sʟ�Fz�*u)k���|G�&d�F�-�� �>��˾�m���x��D��E�N�a�Dm>K	�T�����0��UJ��&HUҲ�C1���#�3ƚ26���J�]8�3�-��X�^_6��Ҧ��Y�$_���^u�8�Y7.���c�ݭ(~�gW�T�W<p�Iǌ�������ƍu��7m����4���:̣�!���	e�M?b���^���]%@�܈*ť�
���ag/��.'���nL�K�ц���fi���[gQ�gV�,i����~�PC� �XU�P�OYT��