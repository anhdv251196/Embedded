XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���������gM>d���`�_����&�i�	~pjwL��e��Y��Z�v8��~���#Y���e�à�8.�m�:�5���!�uY�,�5�wQ�0������;�V�O��"���(�{f�֮�|�rH�lc�tހy"�j��kڢ���-��{y%����_�՗���CW9ӥk��9%���!���5�M2d��W�;Hk?���|b���Y��q�Sܱ�#�?$���&����a�=�s3Q
��P;v�3�f��6��팭B��+=�����]���Kw��*�Υ��PǺk�ѷ	f�c�cI�v��Vn������I��R,z�OAO�%9ӱ�����}v���Β�IR��_k�xO!���z�4�(b,F�Rs�7WLupI��Ϊ���Sd���}W����)�	81�z��Q�嚎9g����H�����8L�$
V����q�thU�2pl���Պ�Kk����&i�e�7���1��oR�j�PNݼiQӧ4�쫏�g�9@��
�BY8,(Yox�U:<��E6���)��=����j��<�.��#T���hRK����t+b��ed'�E�y?�L<��'����uk[�,֐܌yi��q��cc�!ػ���S��-�d�c������"J���C&|=���o��5K ty	���ɩq9�U�J^WA�s�HN��+�UY�0�1�PE�*�֗�/ZK`��ӯ�u��ngY
� `cܖ�ݸXlxVHYEB    6fd8     c30㶲9icpy���+�S����Tp�d�$��J�m�ĿeҢ����V=��i�S��k�6)T�];R��t����2R��z��<�۾7HK�M�B�ڀ��l�Y7*)��Q�n5�+b֥�-��y�:��+�U�H��((���{>@}���E$)3#'�=^�i����t�G���m��{��;-�3G���c띉��	�}t�a��Ɇ��JG�'�?�%%�x������r�V��4Y�\�)������0�Rt6�QF�̅N�$�o�Mc���e�6jl��b��-�Sܽ�5�a��)��~�`��T��������W��?k��
��÷*\��L��|D�H�,yN�
'f<��Yqu	C� ������߀��b#6�S9�����7N�� �g�M��V<��N����JII	�BN�pOPu���-�e%��K����y#�-i}0E�`@�`��|��.�)nI����:�T�W�S�w�.(���g��ן��0��%= H`�wJ���`�i���NI����r���XW[�R�u׸��R�9l-�H�:Z��	�G����������Ik`�Z�/���~˓牤�v,����A�b6i���]�v�خ���T��W��Ή�O��z|p��)��Q*%a��bk`�CB�*��H�]���V�R�&/�Jx��Gu�|9�ןo�PJkp���IGc�-$鉛*�$�W[Y���^qS���X�����D�ر��"��L������x�����X~�A+�x&>o��V��5�	?br��d�z$�_~�i{� aU�iB���|��{[�./���V� 3(�,�}�Ӏ���0����@�z���k�����?��Tr�m��\\��!]�͓#�p�`iJ�Ҝ	�6�X���R��VZ�>/�d�r���ߗf�|�WaG�e�>�~�-KU��}��z�zkb�	�Z������
����n���n,{y~g�+�եo���<��,Σ��})�L��h"ܳ�����'�2 A�P"�_@�����	y�G1e��G�co��q�A?�H�����4�2C)8�9$�1�6xpz�Q�ı�Uks�"��H���S�yԣ�37�Yd��!;��S����T&W��?��a(ܲ��ŕF����>�)_�a"�8��f����*��D�P�r�	�*^C�/��f,Q6TG�_r�= �H{:��u@�:�s.Gc���c�?P�6z{���g�U|�d������T� q�uc�-��d���/�Wܦ�\�jw�F��ѣr���i-�8��N�[r�w����'�I͒L��w�	����2{��r�����QuR��8��L]���Q���qHG��7��C��``E�s���wj}'�k��ڱu0t��.=�������n+o�M���D�.#zm�!��-�����vE;�+��Y�B���l�@%@��%�}� ����Z�xǃ&��\�3�À�C?`>k�������T����U<�@_��a��e>�>����渭Ս�^9��%>B���B2�g�9,��W���������j��̣6��s���w&�2xv~lH
��*I���"�V�j�x�5Aϸ�XȦ��41�^��!� n�$��bDR�kz�W������Uo�e�X�17��"�� OI�m�Ι���Թ��%�p��=!�~�ǔ�~S�g��ݐ�YT�,�9�#O�j�~�����w���b������f����PT��Z1���?�f�aY\DJ��WZDS��u�BSg�π{�(��nS�Qf�f�u"R�b`<���sM��8���;]zO:#�8#�i�	��k��;Hy�bI�	���L�w�3�#t����<r�E��M	���͉l�>-(�E%X�d�,邕�G4JV��P	G�M~� AI��)$Za9�G�e� �I:�f�vq���8�T\���ĔK���5�q;6y ~�hԸHp��4�@Y���9s��bk�� �`D=�2�j��I�l���|���)[N�>A�A�w��4?h�ǳ,fK�*X!�����5�7��b��N^�0fc�r#�*�Dap�kc�rzv��ҤhQӓ�	?��	}�Vb�^����Q�>ͻ0����Nb�_�>�?>�����^�ZO��)T<�2����@������oƖR�r�~���A{��J��̪I_:�9�D��� �̾/�p��:z�!���M�M������^��L&U7�"ɦ�N���p� ��,{,�����2 �:�Cչy�����6�Vcُi����:%�"\���V|E�Є��	P�~�=$^��*���M�(�ŃnGb�r~&�+��"�M}�;�s�1�dǒV,U��&l�̄Ŗ���̟�/���2{ܶ��+�q�爞�7~N b/4����cI����NJ.�L���M���u��gB�'�q:��*�����R�V<�
=Sc1��$l�C�'NI�;�|�rg~�,��ɩx�
a� )Pʋ7��T4�!l���2[�Pkڐ�7Y�Z��%�����6ܨ'  3�t���5T7�e1}O�X�� ̿�,tgz�$_��X��P������R�Ϭ��	ūZz-���X��m~yLZ�j`��WS>�g�x�x~��%�&	��I�%�ڟ�.S��k�˅�aDu����>W��ֺ��;��z���][E?JI��M�"�aՕ�&�?�GOE��� �?7�\��/��XF��i��}��]cW����Kc���RQ�?�b^p�M XT�N�ܷ�1�S�b'�������r��v�3�IB����b�L��3���N�4�9���K�Ia�G��+9������i�(�������gͅ��?֫�5=�LH�`[j�z7�q]}����X�]� �)x6�2q����'�t)x�nN�Aqf��;֛0g>M}`q���1|�򎵸5þ�^m�u�^Z� �H��]75�������3~.DHk�S��#{ivB�����&�ys7��$���	b1Y��|&�t�VNN�B0F~��/����J�.��מ��l!L�Z���cdRà�1�E�>����;���cT7���c�l�?�hoOL�f�ꚗ