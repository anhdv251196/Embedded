XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��;O=j�?�7]d˷�K�[�g��A�
M�uW�+�d<gI(�b9���A��&��B_�G�@K،�G*}/�=�VEh�'Wkx�O[��K_"({�_�PA������gV�dDL���:�HR�'B���g���v���-w���<V�	�)͍���������s��'�����߄�$���� ���q�H}��<~�\�sM|���@g�4w��n�pv{��}(ܣ�ݑ���<W7����XAz&�Pւ���X�ŧ��tsZ�\��(�e�*H�i�'��!���1�@�.U���в��-E[�8r4
�H
���9��A�K�M�G~�l���t�!;�J����Ӑ�f���dA����wd*,�]3!��v@ߊ~)��!�Ჲ�2���uW9J��C��n�w���&�|���$d�&ɮ���E���U��t���0a�-Hr3���{
�c?+d���f�r�=�?�zLTcQM�^�Ѧ�l�Al�����Бߵc�:�%��W��-)hb��_�|�#c��c��K+B��_�6�c�d2�S��ȹ;K���E)*��r����Ở�0WW������?AbRk�^w�l5�.��˲c������3d�n�NA�+Ҥ^aC��(�[�p��!����Aޣ�4P�,���#�����L���t sEtp.S�d��]��č���+R�'^���H&��bAE��f��d��H ���~ҔŁ��2�o,�r�-X�;����d��>���XlxVHYEB    fa00    1960�}QƟ�C�y��j� 0c=�O�����q&)3�z^OT<�.�DZ�s,=,b��r�5Ġ���e�G�[qi
�����Pϱ��yG"U����F��n5X� �X$yL%P��H!������4����o�Hw'�9O`{��p_�o��/L�^ �)D[pE��gʻ<I��N�@#a���~���U�	�!4)i?'u��q���y�fTJ������˜�7�G|"z/� �nlRo#,�}f;��"�i�f�T��������������KSL��V���un��׌�ppS�����6����=߬��E�i'w�mUdkƲ"N��V��Nz��a�F��<��[���~#�銦����	l�j#�ߞ	�Č��<�$
�㖷�p4�	ޔZz*�L�bݜ�b��5.?m�GY`�w��۵.Q�,���~2걅���oUHD�Kp�".��~l�Ӥq����'
yGO������,Uhy���K�H=���]{6�9.��͓}	�&]!J��ѧ9�v}m�Ӟ�����d�<v�S�+�dO<�e7�ʙ�P\���jER�LwtF�H�
��?��FH�t2��+��.qz��C�c#��zF�$��*��.rp�E1M��N���Ι�>���	z|��#��Zu�|�B��ڊ�%��C��Kȸ�ہ}
o�6T��_)�-�n}`Ǥ�>�c��|��p�:29�F>}�e�&ivH��Cb�ֹ��G]����B��'>T�*�N�2`��L�gY�y߉����W\�g��+�d͙��=��Eɂ'K_�m;h�O���j�	��D(Ѐ��
��ϛ�<ӽ�Ya'�x�輅�]��:��c�4&������m��TƖ�ʜ|��h�G�u??��E�/1�I)�-����������,~Q������u�ںzf��e`Å���$@��+b۱�yti�N\0Jq�|�0ҭu�[S�}����T�nI���Y4X���&1?��`E����f��"�i��eR�/�j�q槥!� R��e�3y�G���ŠA�I}�>M����&���C7_P�INaL����f�g��/�Rj����5x�%��X�$��C�=����$f\����m(���t"�lN�'S����J�TT(���1+�vN=���W'���6^<����׋��뮰	��b���1�] �g�3i,��@�:��]�w̒x�)$�s��0���<�� ���J!��Ŕ^-G�c?�S�Ҏ�� )L[w�R�;c<3F����ov�Ǩ�`u�f���M�F޳���K{p�NxDN��s��X$;P`Y�n��8ބ�f5f�?�x� H�r]lO�𯕜AX�-+)��F��]0 !pnJ��`�;Jgq�10��'��0���F�2��!l�yX0�%@ [��n�$�L`=�V#��&��u?��Q$$ˎ�W�����|C��U���S�� �+e���1���X��*^�k�^��P4������=�7��)�qRߨ�7꠼�w�)�G��J���as4��g�
��$z�%\�!6&�N@��Ba�.k�*�8,a SwM���X!A^���
X/8TozFʃݿ��Z�|(ՙs�f-"$�Xxݟ�a+m+������Z8�}��JFq$��c��em��S�z{R��١���׊Z��b���T���������sN��w��b��LBۮ�G�Q�X�)5�ǹ,1�-G�ʱ�'b禓����{x��K��B�>��GUvX>6��כ��u�p���(��XE�v@�ϵ�r-���U�J��f_�����1E�_jM9A�P��w�Q�}'��w�s��#'j�w�6x�ו�C7���`}̆��K���E9k�%h�����w�6���E�E�_�aX�رW�a�Nf�(�C��%�Q+3\��?ڇx�B���	<��[��uX����B���&�K:��?�4��L��y>��/]!�R'
O]j�Ѩ�WA�ʐi����t.̴?��Ыx�l�f���ZD&�؁�|��@KL2�yI�&O�;���ul���v�qߛF�et�@F�ϩ��)�ijnmM�\�UC��ߢK��V�&"�K��T� Q��nȹ]�9۸흨xIqCb�1a5&oN�ށ`_C*mb��+��������f�@�`#�H�?���_�:���B�.�c��Zw�W��G'���q�XC��q��Zq�h���C�zm�3x��h��`y�	N5�s��g��� �-̚V���n1?��D� ����V��f�	/1X�����ﯩ���
<�K����:
����B.��*~��J��b#^m��桾��'��s��wDy�o�b�A?<|���GP�5zW_��;ZH��O�lt{!���@�MLd)	ӑ\��T? w'�%������멑*53�aw�~Ȃ��t� Ł%�Z]&��	�����D���?�[�� Ĵ�a ��k��̱d�����i��?yX���㮄-N^\ƺθ�T�Z�ɤ��S��0;cE�4����I+�YH�x��&��˙B�0�/�l������m�sg�9�0hW����n=$)�Wx�.��sVV��}
�aȞ�H�7Sę��.ڗ�qv���0u�X�d�<����4��D��:�Iʋ��n�����.ɣ��/;/W*��L9��6�PP�ldtL.J._œO<���t!�
q9��51+.��ʠ�崜o> @(Ds:�+�3�I�gJk.Epvt�Vk�юt~4A2���Qec�[X@d�j�d)�P�`�O��Wj�ʇ�i��1_��AI��:����&~6�ؐ���%�
�?r�[Aئ��Q�g�dd-J4�ږˢ-�E����BnGS�u�'t(r����Ƚ���~��ׅp��d�3A	�C"��|��������6���6����-X/��6E+ޙ�����%�qc����h���2��1�hؙ��Y6���2 d�o�3K���!�ſ��]�qW^�A'	�
���g�|�����s��K�@���U�T.�OAb�;<A2
�\��S��ًm���[��ll�����(e�@ΔS��DN���:X��]D������R?��K[�|Һ��p{�V�\s�^;�Z��]���-\��c�ڹ�����[��}�aP���c[t��N=�V����II!�n�[/#G��Ԉ�ƀ��&���\R�Z����>��y(�h0#X���x	�d�¬1�W���R�J��.��Z��f��􇈄
�^��s��L��Xxz�P���x��%D!�-��#M$��^���-�_�"h\m�MM4v����>E� uoc�؋���#8�h���n�&��7U�����޽����4������;����GH�(�^��"m\�ڂ�ă�l,���d_;�r�N�JL�D�S0��P�9S5�J�׉Q��.G�x��� �'ӹ�Ĥ��������ZL�{�9�m@���°��#4�b�JE� ���T�_� ��4��F����J?1�\,ԍѯevk�N��M����/�EUA��r�|w��o�h���'c�Ϻ��4�r���b�n%���EoEw����j�M�̞���#w�Y����Ԅ�b����}��M;*HngƋ��(���J����DN�E�1\LZ����H��n���7T��UtG�7Gbm��#ň�ڡ���F#���x��DԻgUh���������D{���(�2y�|{N�I�
�� �EJ�"ƴ;(�F� 2��5����&��o�uB�ު[n��7���BA�a�{o�ɨ>Q�v�H��oOԜ:�dFw�|�%��s�a~�?�����W[��2FyU��́F(�&%X��IާtP�xD*icB��B���%��@�yJZȩl�9�e��6���� oɬ��]�:���!p��2�NK%�!a�񌘵`4�@ϵ���X/�P;�m�(�D��)�˞��F��1I'g�;f�Bo����l �Z�o_�q��-�j�a�#H���xZ��T�̃Y� �诳��jY��s�����<-��z��Q9{.�I�9��&���7j��wZ�b��I�w�z2FU���l��D%A"���C�A�m~k���	��ʒ���a�!y�H�:P��4Gƕ�����ǡM�HU�n�R^&r抢��6O����r)����1m!TA��Z��A�̩�Er�*��j&���R�肞��-�5Ы�b�ˇ�<:����S�t)�$n���˘���Tc��$аZ�lt���{X��7�ve�ܩU�e���B���.�ڿ�F�	8%���-�^���S��E�(�͚|=%�w'�!:��[Ԉ��3���X5 8�U˪Ө�t��Xms��F�Sa�Z�Q��Q
��DU��m��Yƾl�t��W��1���tO���'�ql�=����χ�s��:K0NE�M�=XU"s��me��Ճ&6�]�K���c������ʿ���+ǣwUZ��Z�-��GyZ*��`���dc�~L���wW�U2G2���_H�.Q��V��������?������=	�N��t�\� �0:{����ӚH+P#���G����K�$b����`N(��y�����n'ҿx5v�#�}��)�Zo� �t\a��0�p>�݇��O��<�`̫��9��ǭ|UNW�c3�t~�m6|e$DO�����"ƥL�Q��Y�uL��k�M�j�����ϔ��
Vӟ00��HJ9�@hnn|�ye�NO h��D�?��E���8�tN����*Z��SU��5�+�W���I����EWN+ht<������z;����̣�� MJ���4�t�<��v�@t}����V�K���g�(b���Ǻ�!��K{	g]w�������η�S uvd� .*�� x^M'&5)Z#�����m'�74��������|��i�ˉ*�	���͞PG���T�'�Q�R�+햍�9��.vm�2�6�6�c��:H�o���,�N�����]�+^�1C���W�2�?%W'N�.��2����"̠�#_�6l���:04/k _�w]a�?!y�#�R�`<�����<bR�?[�p�T�Z�(��� ��f�[G���E�/&�I���nJ�;�4�,���~���]f	���G¸��ID�A��@|�Mc��u��rgր|j��o�
[�hz���*ڨ�>G ��q�=2N��
pF60"'�-�:�z�ZZt��0+��(�����`��t,F9_�=��W��TO�(��� @[y�a�3(��+FE��7M߇���:8]�/m�a�$)x��p�����J�]؛�e�����5��g�f�L�>r�e8�ঙ��A�&7K<xrk	U���E�@ؿ������pqjֽQ��z��$�,�a��m��~�D2�����؍��r?�����_��7�)'�ϼ���4-��X�>���NY,n���4<�G��6L�S|M˥L�ⷒ�~�<	}.�ɧ���,#���(����YR2_h}j���]�d��8�����������	���8�C���ʁ���������z�g�P����H��_���`y�'/P�U��I���0����5�^�<�H��~A�����B�2N�@L;�6Y��cfP
np�ӫs�f��u48Q���;KV����pY�엏#�k�C���-
4��I���l\�ް�CJ��ո}�*�� �!\�	����S`:
�����C9i����;ung�YÖTd
��k$g�8L��E��>q��_E�C�	��(5 �l��b�����m�􇡎��1�n}.�*k����MWX5B��S�*c�	�˛�C5|���/DV�B�	�ީ���{�{ߐj"��5�c�{�m۱�,�ꉊQ�ĲV�e�ڸJ6r��:��IE�J�i;d`J�.Fr>��8�P�F���<"��a���#;�Ë4I�U��+:"�*�IrEy�&Ǹ{0�'��_�=c��\c�t#��z�.)Vsͽ���W��N�ǆ�ŀ2����ҡq�>"a
S����^�:�I2R��j�E���|��酹l�"��q�#Tn�������6�Ε��ͅ3	=Vz:��8�v��{�W�A�����lƌ�[R[n�j�U�I+j�o㬑��yV�X�	*��p)kT�����c�}�E�0��>
J?uȟ��R��(�� x���j'��̌���>ʖ��n���
�D��dxSȯ"U�� ������������ "��^h�?	�J`��\�N|.�,^����^��]v�7�X_�q�d �
=����5��������1�R�u���m��"͢i���FI:#=ck���M*��Pd�Ȇ��@X9;9��zc���k������̰������� nj��r��D�V�m�XlxVHYEB    fa00    15b0�01&��G;&���hd�9Id�}���˵n���s���^�����w��a� �,��r˫I�'�f���#"��ttѽE�6�M a*�YB��7Y=r��#����#��?����"q��N�����Rm~�B�P�B��F�jYl!��Uh�"��{A�O�p��t��t�';`��dR���{��tN����Y{�Z(Ó�c�"\��.�&��*��|2t + R��x@8I[R�CY�Q��/d4Y�V;�n" ����@s��pMj�W��v����4�ۓϾG�-*��  �Q�	ըb7��?H����T��ZX�ko:p��{1�YZ6�ز�|(�q-��$&
X@0�66���a���YQ�f�Ǧ@F�S:.�f�����
��_��`�>�+�x!�%akN��R�o�<P�~1�����ǭ�#�@�I��"�7��+m	y9���g�O�vD�F�g���*���Fv=�2'Ʊ�q
�=��5�M�d��gB�op3�F�=�.d��Z�;϶��$"�r��X�+C�o��aX��<�-o�}+�Ґ7�5����W
7����gM]�O��P�w	.���X	t>��}�L{�%��@A�оkxVa���3������:?��6��57 �.p<$T�Q���pW�'�jՃpNjA�^��e��I�1�;U�9�n����9�����h_�H�+���6�Y��:�3����f�g_�q����Z��4<8��;d���1�t��_ �g��Rv).V�T�'��y�<O�����o$�4$XXl���l�ѡ&�f�I�&�3I|��xԇnY�e>�]�]���\
�7���'��O*FѠ)��E�Ш�>��-3���@.��zV̘@�������po_��%U�2-�&
-�X�$�Y�uM�h���rf5l:�m������]���K���&�H;e�@�e���}y-��a}��H�&��}r�t��5K'��`��NV�	�H�DN[�����*��^:��&
�0+i��&2gP��G��q�Hո��*�@�T4-��0p�#\|49}�fD��o1A�oI�$RK�^���`BK��LB��qD'_Y��'�����eN��	��(�NĢ:):tb�&�u}HW��*6��8͟q�$*;J�{�5|� =���{��:��#)��܆Z�y����v���e���M��Q�]m4�z�~=ۥkJ2����L�a�Ȝ�<'��eܑ�<����h�rX"z*߷����������o&���M^�x̆K)��f��2�㡠GŐ+����GVB��WQ��+<���x�4XQ&����[�i�)P�v���˅@�����D>ӂ�h5�k��e����M��8�ǖʜ��e�xA����t�+c�q���F�+fGlߤO�tz�U_�=c6b�ey��d��ǯ�do��ݲ�Q���!���(�����+9�8��8�#��Q"(7���$HRNW�̹*�@�==?Q�u���6|4�e��	f'i��V+���Һ2(;1�0�,̞O�+7�e�����Th�l���V�I�+�t���nڠi��k�,����sdp��p'�w�q6��Z42���g���r.��g���!�n��"/�e�p0���p�UZ$Y�E�O��N��; *"|=2E��]������aB��!�~���#3Wk��*��ܝOɹ`t�(o+���z���W����qܐ�t��Go�7��������Āq�Pp?����l�e��RKO��
���oc�'�w���/VЃ8����V�������-m���d����(����Plكbf�v{��2��:�O M�Ui�1�dG���ܔ>�Ŕ��&�A�a�,b����)U���}K�#����!w�_�������'q�[���9R��v�ZȄ�.��H����=`RĆ�b� ���m��M�9G�(Y5����ms�i�b�,v	R�j�WBA~�qh-��WIO��c�	���c.�b��S��2E�����
�D��������Bh':$TQ�2C�H�ހ %�����J����J�%jh�=LD`� ��4p�࠸��؎/]�o���̑���n����@�^ѦRgƛ��9�Y�j��a��J=�5��$ p!@���������̗���"��77�XH�C{�'�(���[E���D��{�E��4�yы\x?�R�^���H�'��|	�n��j������VC��	Wte��}����IH��e��[��	�dA�Nz� q���y<
�f��E���+���j�4*~5D}#����h�Oi�Y�r��y<�	H'z�<�����M�]�!��ݏ�6'�~�ߠ�E��������8���eh�;����k�Џ�\�>���I��9K[W}tA9n7����8�������p;G'�͠�R��xR$�����Pe���_��'�s��S�2PGnNH��ǜV��N�S��+��h$��@�a��:����.��&H�Ʌ_=�����2z�ZMw³�=�Ϗ]U��ŔR���m�\��7����:�N:�J}�r���TW�� ~NWF,�a�%_S o�BP��#ݿ�f��N��=�&�ky^A��q&�x�n��p��B*}S8'�~��=�9�����!@�G`CE���\��Ҳ#rk�� <Eʘߴ����2���'kֵ'R�p��юܫzT`�d�hqW�/q�@��#��.ьJAc�nIK
4
�����)!�ǫ��k���~n��2XM����G-��΂�`�XA�[ '���ibtZ�?�3�|T�P�a�۱���f�H�}/��*��,�w���7Wk��߷g��ǔZ����|O���9횋+�3��!�'5[�8�'�Յ���H���%���9������Tea��b0�]R���P��F\�e����C{�FR�5�Uu�]F;�υ����I���XN�z������xby��gA�lUĎ3�f��;��Q��qJ�(d��_u���r=SL�m:��՟%̔��Y���䔛)�ԝ�J����`&b4K	��eFź'xo���`F 9���o8N�&�U����cA^��H�'Ŧ^ ��9�1�k�!/꫷�HQp�24V�]��M\++��+�� ���?�U5��vvf�s8���E�C��O���FCNKγ7��$�R��aWr�Eȝ���rH�3� 2�"�����F�̣?_	�������͌��A�7�}�T���IW���u֌iJ�Bͧ�[��o9A|�!&��iiA0���J���ƠQ�3���䁍�f�ni����.��i��q�ڜɦ�R'
�s��d�Rl)+ۙf��Z�	�l
��DZ���,���L���,���H�tdѬ�V�+)h�t_T���d��k.FJ��t4
�V{B�see��%og��ޮ>�*6Ό�Z��o/�2�_²����y���������y�Y>a&�����D�r�6�w��+�kd�=��
!YU�J��`Э	��@ā����L} �u$�;�������x�y��/��/#�,U73��f�(³R���$��{-���ӝVAQ#����<,{!k�v��SR�N��{��x�[AΛ����$.�H=E5'�k"� ���!�c΅�jy��<uݶnq�R�>����Y��gpY�vj�V�	���%vg6>��jn��1�@Q�r�e�Hhd�E�u
ۥsw�-��8���ݵHcEdڰ�S~���]F��>\�co�DL�������(AUf^"c�R���@�/����]ׁ�~����CMJiN]���Z��Et����^�@Y�֥�X��|�����=�6%�=�9R�=i6.����AH�O&�'&þi��w_�n��*����A��U�
�cFڜ����_�C�����]��~�6��/��{�@�� �x2g{��I�hҭ�b�]�+�8�g���F�nR3k��;��	��Ҙ��/���#4���;g�&E4���Tr��Ty��k6H���ʼ-�r�<�䡯T�b�-����p�@㵃5y�b�Wߝ�Dy1&s��~"(؀/eE�f�y���0!10pi�h�U��|�ـ�DQëZ�����Ș�G�	?o�M�X�p�9�Y�mE#b}�W��~�B��/�͉�-z���t��屮�At�Au��h���]�R�D��Ec۴���%hB������6;	��`�����~恐ā�nm�j_����_���cA�y4L"�T��ǂ?����T�In��g�|ʞ����Զ٬��@\.��)U�CӜ��m��:�|������
�Y[91�[��̯`�	x���9�$H�έ�W6�$9�}���¡�T��ك	�fZ�λ�sh����q�о�U�Ϸ_~x$q=M�6��6ۢ
�'�5"�Y`��WC<�����	D���/�{��TaN
pk3�b��F�RE����=�.I��*��/���y�!��ɢ���㴥�7�kY�\L�Kw5e�m� �4K-�"=�Vdl艈�\5�� ��R�s�"����^��}�8�w����{*3�r���r�/�����.ʬ�HT�#��v�2��ň����N�ȃ/������=&���@}i���)x�)p]��q}�Үr@��,����c��A P~�w���r�w��16d.>
zx���L�zx�]�.]=�8�MFr����N5�rj�/��6�b���<���k.(Fe]s��,Z�ۭ+�)���b���?�~kJ4�5)�.bޫO÷ked1v���+��n����!]� Ai�N�Ƙ�c�9�@�*�	�-�L=hL��g�L���օ��KA�f��6x�F��(�4F�
�^���i�f鏀n��kݎ	�xU�Q�������gA���,#�r#G���X��}�"fU��:h����^�$�>_Zd
�%q�ʔ����Q����ޥ.�n�Ś�i�ǝ�\������W��bS��Q������y�)��l���}�wċ�p��7>�$��
Zg���i�a,�9z�俾3=���i�$J�����Y��������#F��&���Gϯ��1����/��@�
�H�
�׮TRy��\�C��7x?���I��`7�X7d��GO��/N�_=5�/�XL*��z��%��غ����|�3=O�2��`v��HpF��6����N1捩�qpO<�[��@0w�ɬ?�]�MUZsqK=vV�,v��C:j��)�����m�g�Cf,ǆ�3=�ww�Uq�K��a�'�qɋ��?"���>jX_�8�.��S*���HP���b��yw�S���:���G��6c�ޞ��x蠮��1�"I�t|H��>����b�ױJ�޿�Y?��+-CYp3O�[۵�v�߲ݙ�U��;R��ʊp�:@)P7�G��������<��AY�~���)�ݒ��&㞳K��+6䞀v�3I�XlxVHYEB    fa00    1600f[K#
�դ&�
� C�#V������sP�_��+�)�7�ᛗa l��adT^v�.Oˀ��A���ʋ�"uH9�Tw'z��\a��s
��m}�a8����L\�P�B�s;��["�,��(�2�Z��hh�7�	ȯ��D��g��o�7eH{1h�ˉÒ�^�	�:<�.Q�[���������&����-k,�1Z9��qF�Ma�>2O�Ŝ�u��P}��W/#�X!���L�	�\����S������FN&�ɴ���ۛ��o�i��e�|��:���&
Nn���rG�9$���HS��#+�_������E��#��'����B� ��h}�D2����N�@e�h��X ;�����č����@hL����*��6�o�=ޠ_e�t�)��dE|]D�\��#?7�*���|M)��h��ʠ^�<l6�ƕ�F��@���ʾ��*�'[�N[��|0��~�����m�<�AM���d���b2��$�sy�X'�}��j��Z�j�5�_p#jה��l��vG��M]�k վ��2R9��F1R��ώ*��0?�8��y�Ͷ�n��?�& ��(���V�R|�g��ۼAċ�,����I2�7;tI:LY�<rr_�v�^��������F����$H�Mm�]5� �%�i�[BA�#�LGp1�u�=�m�n
�d�\4M:����'ZÃt	���K3ߙ݃�=I�� V�i�K>>���wIۺ��10��� ����O�/8A�-	i��w���c)�i6�{>�Ϲˤ'�d�?��.�8w���+�z� _�x���e��>_����z,|^�}�� +����e���|�Q��l ��m��3V�Y&��Ǌ�:ϯ}W��� �u�~�F� ���s���olI��ϐ�-�3x|�n���6G�)DTķ���!T��L�D��;��Al�]��?mh�*�'o<���N�x�&\
 Ҧ(n5����͔D�2ݎ��nKy�<�K����0���AuC�Ѷ�j#G�j�}� �b0��7���c���Rf�#�`w��hp!"�-�+B?�Ga��v�������>�) ��8�2Z�;圐�֫%/��I2mpvq�޻�Z�ix)�TG�{�b�����e�%�T�^nH�>�Ks� �)|�(o�NkcA��y�;k9r��Ѕ��:�m-�%�����lM��)�Y[�jĬ׏��GV靸ᰨ���fr��[J�1Ts�e�Ml�-���O�J�J�,pp��Ũ.��I�4�g�Vmr6�{�
b���"��*@]�����7z���5�P��Ak�wc�����#�~����)R�s�Ę3�%�.h�Y����W����uN�-y�Z+u��f㴃����m0,�����9��ރ����ouF��4w�!���4L}\��w�:�,�-����Ck��.�������8���H�m���BTLW`�wtv�����(x�.�v1{�?��#R	Y�]o!��8��$����F~����_�n ��ҤR�7mfE�R�"�QMPݠN-������fp^��gόf@�����:����	�-�;��E95`���WQ�Y��Ҹ?b6��Az1��(�%�ު't��W�'ȣ�V����	�S靆ڟը���gK G���%S�<�I.�A��=�ټb����B� ��ɩ���)Bbh���t%�=R�v��#��0N��tb>�O٨� RzɅ�2L���� ��7w�u,�-��4U%�O�Fݽ���-�ɱ��gʣ���6�z��Y#�0�0S�6[�� 3�и#\��#?z���hX�ꮙ��-�L�=�����댓��U����n����kg�Slgp�> ���*����~ ���7�V1�Ǟ��3ب9׋a�t�V�~�G�"����N=޸����
���P��[��jj;�C�,���U��0u�
5����]?����"��ǖ��[ɤ�i��~�O�]\�4Zm�n5TE*knE<��yG�U����� ����^"U.|π��u\����T�	��I�8M}�iJ�-n�Z��5��%�oG�@X���w�ޛ<���n����d���=���yNe�;�D��RgL7Nh��o���X��)%�����U'��Ң��> �F�7 Y��c����<����2�Z7�pwH�(����T~wbg��S}�M�G	'C�������	%� �l�z�������߁��Ά3��6�hw��5�+�\��d�W����El�\�ϗ���$x�\s�.��iLo�z��
��FK��{ea��:&�'̹ٝ܈K�0�?>N
;!�n�̧7Ŀ��҂,|�S)�JCR��v=�	���$
��<�]B�ַۼ˅��4��ރ&J�g>�
�|V���C<�O��:mn'���6���+-2־���l\ !��ڴ_��]!�|��mxH�����Nih�JVhZeoW��Q�%����g����Y��������)�v��9bu�>8���`�Ә�& +�`s$ �b�<�����A5�"�C/�bŁݺO+�dA1
G|�9�Q䙣O}��)"�D���fH�	Oo�������2�l�8T�ڗ�r�Ӝ�QS�{u��(>U.DQ�:`#��'V��ìr�S�O�*D�����c�use(�g4#��7D_q��Q���+	�+���T�-�?C��t�?��&�7w�����6�4������8 �i���JΠK�1������F*����'���{��S���W��H�V�n9������Z&M�#X���gs�Õ�E	n js�&��G�¦����f}k���S\��u�HД�A�Zs���s��k@y7k��7!N�)��Ā J{�w����9��}l)M���"�����i3(��<��a�BX�ؤ8�Y:.YS�D���Bݢ�+g��[K�X�ysd�F��v!���B2���Z2�p���
pO�z�X��*�1dM�]\ӑZUҬTdV�^�+�sO�:6LwK��.��^s3�|GjQ�p7c_C�_~��q��2m�@"Gw�J��y�u�1 ?��}���2Jr�_�r��|pPor�-����X��Q�`�|L�p�
h����Q���T��'}󹣆B2�����$+���� �� =�l��kS>z��ܻ��paӼz�N�_9��zQMˎ7�i;�띱%���m���~��'�r3oY�/k�����$��,%�b^ɵ�L#{7m��]�tb-{[��̾�O���ӟm���3H.کZ��E-0qM�b/f��4�����-f� z��s�f�pKč@�d$Vy�~��?O|��d��K%�+qdp��������}v�
��G�ҝQ�G�&7�tX���Y?��Ӭ
�-$���n��p�g�G��E�;vsþi�TK&P�8��!W�S��U��?4�%.���K;��3
|x#a{�o��w0���s��6���
��l���U�T u��)m|������%'A��d���t���{w	��鲦N�5�f���џ~����I��ŏ�1b��m��څ��L�Z�ɚ&�ۺ��������ȳ��h��l��t���3c�ǠE���v5�Zr*l������'!�-__E�6��kD0s+bƄ{���e-U@��m���^^*�S��8��J�&{&�B4����?�Ƙ�cbT�V?SIn_s{{;��O�?%(� �\����&�v�?�� a�vq�n���(?�(h�/�>�
o8������v�U1=�~��R����P�#����ɽ�"'Ɖ1�'�US+ۓ�&�S���5B���Τukߧ�W�]�p9
��C$�-��(��{o;;+�݌ge��jvZ�XL�K+e��<��\&�2�>�β.gG nZq��B~�Qq�l4��=J��dj�-݈��g�6<�H�c��#�>�<&@�������T@�!�풷�����5(�(�8N�۹+�r:`͙�w*"d�z,!��y��w���̕�B!�3�	2/�A��E�\9�f�_�8�M�׌v u����pAe	r���]Ʌm�P��g��bd}L�[�~Bs�	��>%�vb��>h��A	����F��\�SΨ���	�� E�!A]8�id�Yz�M���e魅�g$7䍨|��x�P%M���+-qDUʛ�1����J}?ӧ'�E�"��@�|�{�I��%i�0v���j_�wg���j�mu�;n�^�&�p[*�����`�?1�m�J)�q֊���M��M�ߺo.ӽ��'28{U"4�� ՟+r �FJ-s�5F�m��H�����#�":��i�r�W5D�79���=c�R}���1����1��F� �j~_w�@,�N�,*m��BY���w��!�w�A&S��F��ݺ&�Y"	��EY��t�*S{�ѳq��۰���w[��y,C^ �oB����\XM��_����E[\Ӓ�i��f7څ�4U�b3��7I%{��
ss��c�er���6|�`�8��r͠�����բ/�I)k�hC�[���Q.R<��*�գI�ł��Ƨ��R��.ǌtw����G�������-ğZæ�珃NF>B�,^�ZY����F��'��U�`���+?���;䝪�,t���	$lE'��c�z�)�%f߾��Se��u�[d��H;	�G��`"@��r�*I����86�Ȣ�}Q�_1V(��Ȣ����&9�x����Ӧbd=^������n���s]?�i�a��ӱ�1��B�.���`X��F� �g%�V��U<�~�$�J�����8�j�zO2��x�T��(�!�),��E_���2�i "LD��r�[.��)m Z'����b�ié���n)����<&�/<��C���)�ƱЎL�^9��`��
�DRmU�R봢�U�x�;y�/	���זS��*�P�upu��LOk2xo�� `���f�C�˵����hIi>f�'�F�9b����Sp���sC_���U-�{oՏ�f�AQ�²���13n��^��N(=WZ�B�q�ɫ�KH����\�ԛ]����������6¯2�m_���.�Q�6��G���,���ߧ�Ǣ��|-_x��A����=<V����BYޘ���yAݜ��Q&R$��@�de�3CO1X�#��*[��]��/$�q�6���%[!i��p���|��!aį��߈�?M�*�<�e��k
og߈d����z������'8��|VP�:�X(-�6�'#�M���+�8V�v��:�ӟS�3�Bsa�FƳ�����5�����*�81�F�<�|Ӊ:$E㣯
�.��Zѧ:$�J$��{�1>���R^��` ���Xm���/���t24_�l�U�oļQV�1o�L�b��`G¸n���� B���-���	n�&�7�z���nFѹ�w?�?d`����1K:|�� c|�i���G��/��D�o@�<���^g	*s\�/��;�6�z���������|q?u��bG�O-1XlxVHYEB    fa00    1630Gw��+�Zy�a�}7{eG�ini�>�/�h�M���Iq��0�n=��R�XJ�Z�j���g��v�>B����hAf��U9� ��+�)�}9�-LQ� y�#H�7���T�R1��kN��t�ώ�U ��{a٪C\Ɯ���g ^�l�P�-r2�3;��T�{�LC�B߷?$����^\,<&-�׶W�5��"�)ǚ-55ֽ�-zx��PY���%.(!�u�i�l�b���G��G�L?C��1�:�z��ݜ��^:�āzD���;#} �(ӌ����"G�8��{�����m�3�����5wEl�8#t���㲻H��j���(�-�@-�QC�1���DF�n�l���|x�,l[ާ~�'h�o|9T��^��F/�������{%�61���*�Ci�D}�D�{�
�Ʊ��� �(W�w�9�j�z����M�c���L��Ə�wL�"���-Ύ��5P�&�rͰ�ˉH�2n�s��W��(��c��ܧ�7�7F��N��7�r�n�8,��nlк�ۇ�������)��3�����|g�QS?�Pe�."�M��0�܎?�MF�nM��d���:�vP��վ���L��1p�f|�h�yPBlS�^CeR	�ϓ�?0 �O�/��\�iFd/���ca^�C-�?����U?���B��i�æ�-��Ť�e��R�]�p�K�ù�);�4j:��~2���C*BY�v_H������u�&ZpVr8ŏ����T]�0GcZ�M�� He��F7�5(QҤ��5�i�gQ�1#q��N[r��n��Qi(铁��~~�x����;�c�oM"L�c�%��d��1���/���Rݞ�3'�Oe�۽�I�γ��L�o��}��&�z'�2���В���֕�N�Q-�T���L��gI�+-��Z��gOEr�H�ks]���+:��o�4�m�؛̼2�oLZ���Iף�s��(2�j�Ovz���+e�VY(l��}��}'�W0ljJ�Б�����@��0�3lf��<}͞�#ff]@`��h`���K
��T9{<^����+�MY�!����ފS���Ӆ���i�!�GUH�薬g��,D.�l�3�J:q�-*c0�P��?A���̗�!�#�T�|��>��i�?��m���?w ��	\㩄���p)5h}h.��9��\�~)9b�BCJ���#��<��٢̙crn���x&�M��k�ǃgz�s:`'�5,��l�mIz��$Cm/׾��Bət��F.f0�9�3�8M5��E�9�ڌ6d�8|�1p�(EV�d�Y��^M�����
.��i�C�2qp}G����%�e�5A�{���d���>��O��B�5q;@��k�Zb�u1�孅��*�r�3I_�F#�:[D��k�Ͱ�6�t�eN�-Q�2v��Mi�?�4�N���ޝ�V]���32]\%�Fd��1�nF9\�؄�f��}宋�)�"�%�Zh)x0��̛�vX^�В>���h��-`�,���Z.�3̲)��i8՗v�`�s�dl����9z��A?uƘ�)���A�%!��B����n��T�Ë��c9�L(���u�����ךGc\�5���:T|����&'�t8zh4ߵJ�%D�?�-�N�[�}'���d�1�lQf�*��U�!����q^��l�\�U3��^��AL�ȿ��<�Ғ��ˈm����F��j�v��+�M��W����W߲���܆q���rGΊ������Jg��,}�R��!���9��҄;��|�+X�g���Mջ�L6�!��������W�#`���!+cI�Y���E���}����ym��p�`����LT����}��Π4l�ND��A%n����� I��Z/qqӲ�Bd�)��� -�����*�d;S����r�N��W}_� PӦm.�qJ3��e���9j����2sq=`S���`���Ι�!���1	�u 6�� �Y(q,Viu��=��[VQ2��Z8�I�m���ʽX��Sݨ����Ȩ��-_-�L�� �җ�ܯX�[�E��NĆ/0��FS���&A��6͔������9��X��6|~��'��X��6��ҷl�� tD��x�C�s8&Yx;yP���{M��~m|��_��3r���!��L�^�dp� ���Qʰ�4���Jl|���]ȯ$�ɐ�x˰g��M4O���4bt�~M�v�ձ�o����[A*3�`��W�Mte�p��aRSHTaG��Ǟ��Ȋ�Qp�}c(�^5���p���p�����s���ƛG|����#��Nb�\_`�5|��� �������>Ƭc/BS�E��(���)5θ���7���\�wT�@|�o���\q���q$鶋:���GI�A���ّ>�dZ�:�꡻"H���mxOb<5�?� p�Ʈ�r��{̤�@��|���bbY���̈/��}�>�i�&F���_�bjf�m�2�xHx�G�=�n�Mb�E0�T�����.��	?�8�����|����-����7��AF�C� P�z�¡����DL������ݧ�"(�ć��Ŧ����Lv$�i�C@�J�H#rZ�A�����R놭��`sQ��d�ď`�OtHK�O~��9�^��o9�GXS 6q'+(A!.#�X��sxx4`DL�ԠtZ@��i����V��X#��K�^�)���dy\����F�hD��_&����6�)�m<j�smNf����q̧E�T�������uZI�ڰ��n{�V�j�+hj��N�,��n�C7����s���*S�����H�I��s�D�ż��r��2d��M��eYi4�W_�7�d¢�2��o�k�T0����R#$@i�$��D�&V��;-G��j�R����`����Ta:��Ó�)s��B2�G�Ho
�0�^���U��y��Qrc=���$�p� Y/��9ՎP�X! ��0>h���%{��e|2��_;�
��2s�
E��0��V�ើ��@�*�4$�=t�b!�q�8@�r�3�R��W�(��q��G�����Z�E{}�\�
aG����4~ʺ[7{�<f&��Z���	�b�*wf@�i4W����oI1S�`�Z���Oy�=�S�����Ջ��P�!��3�Kؽ���4{�^�U�kum�2�����o3��h-�ʆ��0}gu&�^ J3�4�`�@)h���v3U�J<�1�?��ҨM�{�û�G(Y��E��	ߙbv�;ruF�·>u;���z���#�=��C�1��3�A�^�H�"?�Q�(���:<�����h>�1�a��8~��B-��X��~�}v<�2��=�v�͎�5}�6?mqlW^j�)5�+��/�[񦷵�W^O8�L�/ֱ������Y�z*�J�O!EK4��C
8�
��y]�>/#;��t�Q[ܗ��6�Yp�1�.�7֡��(5"W]�R��>{�l���R{)�3>�_1�:]ru l$��;�b��j�2��^������D�ڸ��`��h�|����2���f�{=� �:@n�̉���GvQ2j-**K݀��y��ﶋ¦_���ӟ���|�+��:�ū|��c�`�Foj+�bOR���!y��qw�&t?�b���z��S���3k�AQ�ʇ�qE���d0��.R[q���z���|t�V��g����I���1OO�5��b�|�D�n�9F[U�o�.��b�үGw�20���Fx�T��G𽸇ȦU�:��K%]�A[���;G�72b�p��5QQO�����d����|�Gq�F�|�E4��yu)�h{l\�	���:�*�@<�.ꝫZ��W�	!	<�imtK	S�_�Up�2���� 8�y��Ѓ�S�CxC(��8����n�j���D �Q\�Q}yI	�];�R�Q�R����AZ �,���`\��v�d) �9(�:����<4�S�$dY����L&f�=�F�>�����e6�
*/Ui�ܚno$��Ƴ��J{	5��O�x޹I�����SRݬ��]oCS�����	
�P�>g`�+��r�w� �Y[\N	��	����ISCαC�{/]�/����4�P�⍦�e�g��HGl#r�:��4�=7u<u�R�t����'j�}\
��M�c� ��K'���@�e �};BK�O�\��0�k�4��s�t�Y�	{�;���U�>O��������G�������M�ǧ0�e��mfg�Ө�+���W�"��w�������	S�x�� O�'�U�tq
�������)a�$�0�)C|Π�.�̓e�	q׬r1ۧsJ����
xõ�%������O�!�m����L��u���.�X_e�ɐ�:&淆��D��VZH�7�By�P6w���p)ЭU��wE�@^�^�јR�_<�֌���G��D���g(��w�*�aY��r&��Cp2�����+���K�ݫ�@���ۧ�܌���i���m��T���]��#+OYW_Ba��v�o�q|B��qo_=��j8L���,��1��KF�P��jt�����(��f{�xp��8�<�I��n �`{�OJ�_6 ')a 6w�)�2������� S�Բ��5;��^f+���ܘ�r�TW�/�DC[�z��kZ�>���ċ�*p�\٨R�ꆝ/�Ϧ�OC=s��rN���"���,Y:mr�����|����!)@��y�A,`���G�]/�FD~-٢aq�� ��0ݴ:�������^J j��E9PQ"i�K��r�?�r6A%hBV�r��R0&}�
3�D��ڇi����Gp��k�:$ܸv�z=� y�|$�|�����y��K�w��Od_�k��o*�{�U�*:���i��
_a�ؚz���s�M)�;`�6��N{�L����qܶS^V���{�2%BO��"�,�b����e��n $�n��|���Mh�������q�c=��cyy�%�=0Z �M9.�o�'�Scrļ֬Χ���h=��R��f��[~U[V渙4І<=��D������Nc�"����B=鑒ݣ���v��]jdeD#�Nvjh��ˑ[d'��.E}�w��o�0�B���b�.��	�\���ē�Y}TF^D�������EQ�G|��$�#��'?-��9˄E�NeK2���4�.v�kX�T�H!����C�|B�$N�����J�ũ\����tCm�Ÿ>��L�?@P��U��~��C��@_G�I �_��U�LAq^�����RO��,�#x���>�^h����$$�٤S��ƗȈ��k�_*��W��՝�M�1����{����yn�gD}�K{[�0�~�~w�1�eu(�uhs̹�����$4H�zA�$��*"@�Gb�f�v�oR������r�CJL�=lD�Ij�.��XU�����@�!/�_o��h̈́`fϻ�e#�1�n�E�tp
Be&�8��1[T��#�Zt�'��)�&����� P;�"4���e�]�Y�>l �V�Y�����?������}8ڥ�%�dT�8q���\�a�eI��i͹�7�W��M&b�I]clXlxVHYEB    fa00    1620���Y�}�����'�@]�MIY4H$����!{��*�ӓYeWm�c�=�4#�s/
-pG��`�ɖWri'��s����R1;��@�J���7j?~<(w���|��7*H/IE����'�y���;Ta���.v����vB�2��<?��o �bSd5C��f1��~g�i?NA��ѐ��Cj��0$�����_��i�*M����OA&%��Kȗ�o
�Vj��5Dv�|K�(��	?e�K����	ú�:mv���0w����a��yZ�*��v5Xh���c�xl=�z"��s`�d�A�!��R�t�n<Xd�z=V�6:���9�j�B�����`��������S�kgŋC58��qajg@�z���!Dэ�D�DD�D��4�y8(�,�Q��(\Up�N��.�g�3��� ��yaW�#�hNJ����P�>�J [������ݟ��1?�]���[��D���A)��O��p@)��sj��%Z�|��o�2t,��K��ҵo�@&��G��6� ���hh(-.B��Ǐ��L�U���FO�%8Lm'Jm �7�T����:u��t6�۵�����M�Qsc�,��T"�E��b�I�N�!��]�� ʱt~Lkc�sA�Q?����C��3��ԩ��VL3Pr���*���=�7�!� {F�%��(nq>�=R�&
?�g�H��ou�^���1��_^d�71��%K��f���3��<	A�V5�Ak���1��C�c�-z������:xW��	�ǯ��H�Ѐ�_U4~����A��C1=G%'[<�qg=�׾x,�n@��i�,�x ^s�n��*81b�A���>`G��O��:���,H/� p) �p�]O�R��]P�٣@2�fo�f�Iݾ��=o�x%��L%/b�ٸ�B���vp���Hm>��D���o
a;6~O�o���6b��U���{�{!?�R�/^ �^��h��Iy6�&[��J$�:�K~�gG��(��g�R�����Qp�Œg0���A�v*��8tB�@�M��{K�;�~%,f��'���n��R�/�#������J���;P¿4܃��}j��ݶ�8�Z��:����sް
�%o�~e�e�����ҭ5�$���_Ɉ9s�꤇�.7��	��}�z;L~Rő�-J�S��j��#���3α��J�ix'�^g��з�N�.��ݛzN�9(�br�=�F�<:[[�RV�<�'OS�{�W���m��id;�#jvWK_��yn&}*G2��R�Lg�@u���h��s"�哘U�<�4LP�Eh1>��i����n�קj)}5���3 ��k�	��*�� <s<Q�`�0���9/v�)�����F��[[��f��uD|M��<ĭmK�~|-8�Ct�C}�nJ�+7���$!@����S��H]惓��'��aQ�����:5� ��7�כ(�q6u��d�
�ց�A
sC�Wb�<�V��w�3���G��mot�s�dcO�<��b�Y�V��(*�Zd��q5C|�C�]3��tʾ��i��r�ObD���� ���FJ+��ة6��� �N�����y�Ӈ�����S1��&�=H��I0or�����rɼ!��\RPΈUeJ���S��C'}j�wv��{��!4���Nn�E-V �K�CV�� QE�c�]�dz�f�V�^w�����1�9Idf�[�b�'Q�߳9_^�=v�+[T����(���zW�DNۗҘ^�:���<.x���ʻ��^4f���i�{i?�v�,�������hc���k�v��A�`h�����ٶ�)��ŶlbM�}� q0��P�)90�n�[��+0��!J�������5m/S�ɐqb�5|��?�+l�t:�1r��͘��@�Hs"%�i�s2Z%.^B�z����1Ʊ���XP_5c!1SkS@��{κE�]�d5���bI��X�&��a�(�ӿ� 'E�IB��L�e�^=�v�q+#b��܅ Ψ���2W����X�������Y�,W�?���v5t�L��������AK[<n�vʶB	���`�� ��ӻ��G� ���.�]����*���TO�ca;W͒�������*/���p؀��>fr��Wy^vh�(�R���$���u�@K&�S��͕��/���/�*,�vb�g֗~��m�zm�a<��}),ON��q���z����Qp<��� .�I�����o�����d��[%����֜=;`K�h�i]�����~�n8�x���io�TiB����`sb�q	�iץ���}�QFr��tb*ϧ�I�R��ͭtÿ�}X�X)r�I����L��h5��Ūl�OQ+�-5�<(.��e	�8�4,�\�|���,$4r����B줴�f���u��պ�Z�^6�;YL7F�k�{�'\��k�;&�X�ҡ=h'�3��1���/6��b*��@�����,VN�hi���6Z||�T��O0m�2~r���z����sh���=o�����%����Ie����S�T�4U�L�')�T��֠�QŮ��\LE�\��LE���B���;���a�uA���Z@3����A|����YL�p�,ICy�����BP�	��-����v�^\NI�4����.,B,� IRX�C`�9^����x�=�q�{a
@Y�F�2n��"=�e����c}Q!�$4�ڧ��e�5EĬ������-z=:��ȽU�e۬t����l��a�j�a6�X�ڟ�%�m�_n�� �Z�e�/w:e�ʅ��3T����X|뻲e�ؑ**��)�D�X2Ҝ����if����8��w�Z �)` �� $��s(�fn�w���,|A��6�s���ߏ�?�)���>�\�R+���3�[v``R��hY��m*�go��)��].���ѯ2Jx�R�km�i?�4.�-��ȍ�	03Mn�	~�w�T�$��N�'�C�-�Z�x
�-	��5������Z�� ��d?�ۘC�KaǳwT�j��X�e2h��Z��]�K�L��p�R^��Ή��)"�ğ� L��E�eBYB
[P���$V�m����U�"��'F�����}�)O�f�š\K�76�ן�e��c|�u�'h�"{���e]��u���_�<���SCm!�X�vX|�r���Y�r��A%-Ȁ�t��y@���I:B���ZF(Ym~�8Sԍ�ҭ�+Z�;OU) ���z
��C������L=��+b���9N>�2�SC���K����Jk2�V4赺t���E�SokXntQ|�"�5����q
~;�m�u�tBt��J���z���5=�jn��������g�aP5ZI���'D�+��%.\ .;��Z�1�O}���*O6z4\�����m�k׳��j�w�G�M-�N�'b��Er$�"�!@�Ot�_?	S��I�J�oX�u����cP�k�-�D�6:�E(ɫ���݄��+[5Vn;��<z�ߵ%����^���(n�d���H]H=@"�%3�t����v�m��u�<=��w/&�гe��$��-D��� �@~�<)�y̕d��a�:ÒJEvBd�/�M��ՀƧ~ϼy�Б��\������a�T��?�덠����N{��?b���D�����E)*���r�n`��Ta��������t�N�<��C����g��mg
쥣���<\�d��<�t��K^�v�C�<����N{�	�����>i�����.�j&��Z��L	բT�{��.�9�
�)�i�`XM,�r{���$Afʶ\��01��+{/�"��7_	�A켸ϸ�XlͰ������:�}>^e���q�+Ж�@�;��;H֒�0��ZLq���C����	=�{^`.�2�r�w�H��"��	[�%����.�h����< �W^aR�V�8�u)F�P ���*��I���)��I�#AYe�e��.��������IϤ}��e��1S��b�?�C�������"g)4럴��l/�a����t>�)��܊����ƅڽ�+!%K�TdTөFC�@p$8u�4t�?���-��>/fH����~�a�JzŤN\@t���ώb��|�e���n.���6�{���B����K�5O+9�F�<�'��'��;�M_՟%P~5�����yK�OE�ҳk#�XU7���J.@�QI��&�	.b�8���aحw�Y4Qkx*�E!�̙���!_>Y��9����+W/��b�9K����&�0�~���=5ڵ�u�Ҕ�Y�盉���+��F���ݫ�9�uMU~�lē�/�S�p���F%ÿP�τ�E����Kϖ�rp�&Qq�x8����{"�����6~T*��$�9p��	���Lz��Y�Um��q��	 M��3^�R�M������úL�)dw-�'.�a��-/�N�y��i�*ru��Qz���y�j�� �|Y��Gt���6�y@#��w�,8��.(�t�U��K�(�i܍V}�ľ�`p��d�I"� �Э�R߷*G8����v90Iqn��G��)2�� �ew%�i�2y���q,��ت9�A�j��3�J��5�j�$�Hs�\=(V�\�Qh
�c[�����G��_����]��q�!�*wcv��]�t�L�W��n�w�$�W��~D�J>.��a�~�^d�8�_��N&,JbHzf�K<4��bl����:\��(l�ld�,��������mw����a=Lf�+���;�Z�Y�A	�]��jh�x=�����i�����̣Fa#�.���4A��[e���|�Zg�_���V,E}�!mIƟ���H��(�
{X����v"IH��f�%�y�?�F��kS7���B��`����M�7�{��A?��1�T�N�n]���5"3c�C��uj��o)�)N��m�����&d�5[�(5S�3֕�n��(�H�P�_c����
ڰx%�@��G�L�m.��O8��Uϵ��ȡ�����3v|ܰ��&��#+jR,��1�*_��@堜���ț0��#RYòr��kiw�
��	]�����a� �l��
'�-�Ű�Иz�7Vb2<H���E[�����o�j�Ct�2�����IS���x�t��#�$�L�:����G��5��o��9��h% {E���� �S�(�e�C�V&̢���/ϴ>ii�J��d��x2����"�!k@�Os�50&�v&e�vd�Q���uU5��[�?uFW��I�{��7!i2Ee~Б�6_�^�����;,���R]����[d��)(�郸R^��C��W�Hig��2�I#<��Ã�]�`3�I6)h�&�;'�I���ഁ���P���T���.�ыs=Xa���\ PΌ^��GҴ�_x����#�m���/pyo�V��)\�\:�#���ʱ�#�>dȎ�_�aF�d�7	[T�&���6_�@��2I����+K�-�����}5�����F��5����.ב�1�����ʯ7aS�*XlxVHYEB    fa00    16303Oyu�u�����l��#�k�hk�P#��ݒ	�FK�e�	
*��j��K;.L۞S�%8��2�|�����L���)q(ތ�]Ƞs�=]4�p�ZH3�,�R�2۠p���D'o%�y[fD�<7M�^b$~H�0A����ر���)����>nH�e�R-���.���`Td\x7�I #�� 	\�{�ܪ8xt'��تZ�f*_���(3fp�`��J1��u&�\�M�?�e*�+�bR4����&�Eq<${º��:�IÌq0��z]�#�5�o��`��%��x'l�(]����&�b�4�5J]y��D�qR��+�}��t#��������׻j��kq�[�Ⱦ�f��ּ:V��f�K��U�m�Kj�E�i�rY�W�ϹȲ>�}Ǆ�+0����T����ȵ��*�w��	����tY�O�H,7���Q��Έ[�DR�~�4>�]M_���2R�L;g\�S�A�E��{�@�5��bu�n͕d�F�#�њ�#������`�),��-Q[�HW��0j4lCّ^�O�G���n��hk%�
���`����MU�3>��9���./jM��6#�#��d[���g��*o`��:�
��* ?��7��j(�5Ċ�Ut�=0�-�L��4*�0�W�}�K��l�S�EO���>8��%o,��a�Z 7k�t[�WcPjz�����|�P܇���g�i��┣��}�3BŁ�ؒ��|a�I;j�<���L"�Xo��� 9��|�	� �e%��\ud��Dh�p�ꅸj�y.���}�G�Z�qAP��M�VҮ�ܬ��V�p]d���j��0}��F���ߙ��τ|����?���2���t8�����{f�=R0s8��`��)����%� /�%��)�:	Y��)��Y��˚�E�@�n_g:M� �u(v���R�Cf�s���� �z�4��	�h3"��Mnh�-@C����C�>�̧���=�B/�Ȃ)Ep: &G�:�Doh�\��C�Þ�.�'�Q��@�������t���3�H����H�9��	'�0�U��;��l�Br��9z��KW,�����w�F�?W^m��qJˈ���}�F.��5s;����2Hn~�N$��+S�Ӿ��_ifd�lU��O�d{���<�QG"�/�Dذ��;�is�N����zl��~�� ����_]y�}n��`1��ݸaI��Ž�syo�,�����􅿿S8�>�c%V���[�jC�-�i�c�g�F�����_z>tO��Y�)ߴeJ� �ә�J�(ڒ,�!��U!��JQ]�r���`�
�*G!�0� �jׇ���4��;� �n�o������Cv�ָs�m�K��G&�U��m�e��o(�;j��3IJn��J�K�^J �p.�4�g�Յ��t9���͆M���۷�7)|g�8��_h�=�G�zQ7�g��?�y^��5��H;�$S�;��~EW�Xx򦨞z���~��`؁��P���
���\"0�Ӽ��`�(b?_ �f��X��')	)`Ľ�ZZ�#�ZǊ���_��%�g	�*8�ɍ��?�-b��X]�f������ !�+r�,�lV5>�}&��9�t�U�u��m�����.0����Np)��?��WA���P�*id� [X�A�ERZ�	oKݔ.ࠑ�IAЗ�K���F&�Tq3R�p��Y_��%����y�MW�@�_���{�$b�|v��Z�wƾۆǠ�Ԓȿר��>�c�@�������p��"&�N���PGe����/��3�Պ9/�����_%�6낙+�>�{x�������k���b�q?&G���ۧF�_��H��r���Xi���`gb���;Z��j�@a�*�5�AGv���=_��!�_AQ��;��`���겵��	��g�����:�^�J�P��0u�w���k{Dv'���|n���~e.%�Jȯ��8�p;�*�,!%�wZ����vF(�A%���4:NSV�Ug=�a�m-f�ޘ��ŵ�~�|k�!�r>�{߹wh�c���B̶�K�{p��n����Ƴ�gب�4�|w>
Y�����=kޥ������N�!أ�Ҕ��S�®d)*��x�f��$���ݲ�W��V����T�5��o{I�t�y���1�R�+o,0x7F���8WK�D�=dKD�^�R�!,�#����Z�6��8���.O���>�!Օ�e�H"����ͼ��K��
���q=�v���X������7~��3"f��!٧��7��?��"��/C���'
R��r�NR��,�hr�~TՁ���l�7v{��dϒtF{���[���
R��7�}�ȸ�K���H���m�e�Vt�+�������|T���;S��8��L������uM7�y��Ø�Mu�Zd�������_�A��d��&	�HL�����evn�NsPP����帖(�� �Ļ��
ټ���+ֺa/h+�V}Ea����������P��pc%��rU��Z����͜�����լ�dPKl�~�k�q��S"-�=��Lk\yE����6B���V��I#G��׀\(���]rd&��)�z��âF��EMt�ሦ���\J��:|F�� e�>缞S�4Y��[ʞԺ˷�#�:TZ�Q���pa�LS�mķp'w����cM�
���������o������o��jk"�h֔�t��}�N�r�������#'L�VI[��F*�7�k�:+1B5������.j��;3��hJ�jI{�jq���I��-�a��\?�����TSM�TE��8�2G��fN"V�f�̨�f	Q��x�1�3�#DP��� S
aԐ��qd���r:K�pNO�p/|���	軪<ޘ(L�l1\��G��&�{*;����ښ?��Win�7��潁�ʧ���QS���VI�c�*�a�(�P@R��d�W����OQ߃"��� �	C��!�c[S��`�B��%��&��OGر����P�������̚���ix���-�5-ݖ��-�A�l���'e��I'�����
p���W͕Uz!�Dפ�_�v�ՙL`_f5@Wyv���� ���͓�"!�FYp��aO/�e��_{_m�rץ�=�uX��U��+*bE���O�x$�?w�J�V�����pU6%H�9�)�� w�:�B�o[L�;����O������W�S�F"�nT5U�����>��>"�a' 'm*﷕��~] ��}{��U<��l�e�JQ��zas�m{�EK�!�ʬ�&y_�Ȕ����u��ϻ��J�q�xP "�}u�]v�b��ڞ�~݉d���n���G$2QGK��ue9_У~sI�;�/�UBU�����P�Z�p ���_ �p~ӵgy�.�����ؤ�� ���c���� �|��u�_���PB�����_`����S	�>�Y�]ƀ$%;�|I�
�|g������ �1�w[��,�h�ܗ�X#��Ã͐úx�D�`�e���A��s�:YS�l��~�fm&	Pz'~�����l�&�L4�w�=Wu�ƣ���=��p�Os�rC�6��B���g���^�Ez5go�����$��J^q�y[/nc�'�{�-��Ң��!��T2#XP˫�&�Љ�@ 7�˻y�i`g;��W�gL8��*��8��w�VG�\�*�iA��@�z�,>W�o���'A��hiQpu��$�s�}B:�u��h�%�ٔ��ȹ���\a%hױ�`b��e�sI��־*�ҹ�pG9:J��`�	ۃ_A�,W��}S���a=P�_@�
��R��~V�y �q3�O��f��/�z��{�1�uU<����c_� ���}������n�������9H��1 �5a��Q�f�7��pkG���m�[�]�&g�D��E����KW$�,�̺*�:O\�2'⭇�6�x��;­��0!2.�2��ϲ�J$�h@��z��*�.���2��tp�x�$_H���آ�Z̍�Ïm��@)���_��p�%�2B�Vsy�vަ��uA���0w,/���{���7kK��]���a����xo� ���zɹug�g��������D����Y�T�o{��qp�m`��a*��ޑ��l~��(��Ul����Q���*��sES�ҁ��pxE�����+NL�?:���������N�.���\㥝�5�d'Z- �ᑮ�l/V�e�/u ��"gZoa���ci�L��($��g���Ѓ����Z+���6*�ͅظ��'c0���[[O*H4�Դ�X�/G��Lq�E$�G���)�](b
�k�3���?�`-KaI�@<h�Ă�>nz�����dr��E� ��9����)"\hu]r���'_�o�ǈ{�]��u>���h9'�/�)J�*Y4~Yo(��zO�MIFs���/�*ϰQ���� ����>�ň��+���q����4%4�3����U�)c����,'�y�wZI7�D�蘒�~}�_k���k-!IZQN��v7�O(�'���%£XJ`uwc�.-�E���{�9��	��r�G�g��[�cV�'�����M�etW����v�b�M��Df��H��Kr(E&J�Lq����2�0��v\�����qP�U�R��\�0PT��:'�`�D�	��
��,(�������?�?��!w��_aʡ��R��韑�a����<��r��w�F��G$�\i�g���s}����L�V�yI����΅�&qӵ=e�V�k[dK0L��dY��Z�>�-���].0<y��n??�N)�Y'���<�!�g��r:�*����gx
r�J�>�'�s8����@�D�~���6���8@ӎ�����ת �g��E��?��`C� %hKƆ�� ���xF_���pc�FNk�,���TZQ4wq��щ4�'p����Y�������טn��%,tD�kq��R;W�|��tc��U�~�h��A��_#��Z�@��e_�����6�F�wV3�f9  ��@j+�mb���|���y]|���0��>��	"���%�{��P�;���X�Sʧ%_��-Pd8R�pR�x�o[w���S2��T!��d�����Ѷ�(ķ����is�q���lZ8@�7�_Sb��B�����:*}[<�~�}�����I�pt���m̶�PR��OV�5	��񪚃��^Z��H�����~�	�4��lR	�jn�>$�V(�.�T�Ř��TK��0�l��H�7�8Ұ����|\�,`6.x���Ex��}%�-h<ұ��=��r��m��F�������x+Y�g�N��F��eΠ�V9D�O������ݡ���?�ۈ��;����yg��(<,�0:}ce�m����"���R �q>=?-�y����T�'�ǩ�q�[Z�@&W���^��K�x�-^�������|�� I�����P��<�4v�m q�I� \6�H:��J�1����ĳ3����UGGɪ:� mb��J�Q�3%j��<��q�;3s6h��ҐCR~VJ��oXlxVHYEB    5a90     850��'9��Y�AΖQ�~#Z1�;b�}�t�W!�:q�#�]7��~�Ly�,ؒq�h��u�f#�P���9w�s3z��Um�3�����F�_�h_+�Ly�Z'�p:rt� +� �W��1�;F"q��R�5"fYe�j�Ӑ1%P�伷7�`Ǻ]V�v�"\�h���|uS��
c�-U�J���,�����s���6-{��դG�e�.m�,ͼ�,�C����8�`E��.��%��7`y����h� U�>ZJ�Um&����I��l�K �X`l��>���<���ý��~j2])L]]ww���o:5��4���;���M4�(?uԳ��b�aU��lg2t$�i[�H���m�W�)5���.#�=�ů��''��0 ���ünY�ߋx�y��J�X��Ĥ�\����\o��C�:�K��ض�~в~��Kԑجʡ�N�j��eF.5��D�ō?4���q�u��@�b�h-�x��'Ή���o�[~�W���5~��/�,S���e^M����<`[X)�7p�|[���9��I,�|G�qs\E��]o栀�w����c��hB��1��A
��]�s�Cc-���KT,$���5�J�l�
����
�#�ҫ&[�E�&�U[A��"b�허�D�op��|)O:ع	�q@1Ry�e;�$�1H�-GODmK�ɤ��5bҳ/bN����\"�;�H�K���"=1܇J���N�����d>��-�>�	Jv��
��x#��v�����\<I��8Ȋ)3 ���P����͒��h��?¯���*�����`u�!�`*��ow;w��.3
��1_W��[0���(�x%S)���	A�^.�%]���#�)Î���6y���M��h��wj�g��,�5c����Fq��~��O��>�b�ة^��o\䇌�S�����Ca�236&U��=W����<m�1����U]�{N  	�i:Y�3��6Y�2s����U�d�ϨJ|����=N1eFp=q'Pf�-�2�FTo	�ذگ�NUWW�}��pV�&��Ig͋�%E�h�	=䩌��1�^A;^Ge?F4�7j�j���% �ކ�Dy�P���Q�$ڿ��:�M�����v��_z��FqN�1�>x	ȸ�L��%oɛ=�$bh����5X�ȳ�(R\�U��n��68��d����"�l@e�;&��,�G�|bK(�~�pp��)蚞������ɒ�QH�j ������o��2Tt�}���ˏ�n��YS�e��$$T@��xX��#� X[[,RU�n~��\a�o_�9Q%��2�~�n)1P�]*��.�������-�;J�7�����|��c�//	����Ť�G��M����V�'L�ʄQ�䋟�91���!�,��?�����Hg)��ũԿ���c��̶������c���;0�� �*���֒����s��жB��n�ehؔ��K�N�"���vKq��P�v�9�E��h4�͚we;m<�^p�^��_ۃK�zfR�f�tq [l������!�*�$����xz��MLO�S���!U��Vf�E��`�mñ}�,����2��e�p�VL��s5R��c�0|�IP3��7�B�M��� _�loV���7�a����7��O
�[�����͒�Sa����r���7�Qޭ�Pd7�`�&Ŭ�f�m���&n�(X��q	�S9*��J����X�Iѽ�0��:L.4*��'s
4��r._㤊Z��D-x'N��D��CģX,lV��9S�_��8�.�m�� �R=X]��|T��V��;�q4�%`��.n�oƐ%Ew�[�fz�u��><�i?/��J�ڿ5�؞I���vn��vŁ�(@?�,���gފa@*�td�JCq4����0����x^d�AA���8^,뿾u0����e	�7ё�!�K���2�CA���t�yI���͡��^��\V�Q�-��(AvUAݎ�s*@�i�s�[�D�'γM��]��~��t�Mt��DڜuCvR�'o�]#Uxб�L��X���G�JӄB&]�� �}�'ǘ��~���v��	