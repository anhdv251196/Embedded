XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���j�NO���}�Z��[���ߪ�D��pX�O8�L~�$�.����b9��H�zO���?�7���~-s�3��k� �_�SuF��aIއ�v�S��r�6H6ʀ��V�,��B�*��A�>�96dA����ȕZ�3=�vX��ⱒӕ+�a.�[�.�|�luP��m�; n����:���m?3��p��f���F�WΈYZ�ڣeT��t_�[Mq2(��T��}A��0}�׍a������;t8zU�U��*�=ǟ�ʪ���i���A��u�+���%G�BŮ�wnb��DQM]�<S�Ol;!�o�0�(��j��]��!�������	�T��W?�ǂ,�v�6�C���i�QXF���2k��9nYa�~�_G�>���ȮU�>�Ӗ77td�fxi&,� ���c�a]�a�/&���B�+6�X����^.�h����C�Z 0�-E#��M)[�`�s|{��Љ'�h�Aܙ A~��[���@]��Cip��Ә�m&7��"�'��@�,�K|�B��B!<�4 ����z x�	��H����;�o�����E�g�=y�ΐ��-
	&x��q��Y���3^��oy�i78��탛NYV't�j�X�����\�Lc�	���׺ �[��>��S��Kata��!�v��f�)�BQb*�"���B=3[�o wj��f Q_��x3�"��_���9P��E��Q��*���"=�-Q�g%��� J�jb��(hH�^��&Ǫ�<1���XlxVHYEB     935     3e0���Ex�$�R#�V��T�˽�/�T{>iO�DE�V���U%��E4��w唯��o/ʰ�����E������_2�0���"c�N�#-�dV#�*�?L������j}�2v����Z�0:#,��]���ޏ��:�'�����M�+�15��� 4J��p"����D�0�qN�lc����(�&�;�Ag^y���ގ��ư��sɜK �w�t;��K��5	9q��5��}|���bp>98B[*H}u�H�t@���ղa&��GC;?Q5�A��+��q���_c��Jq�Cr+�h�aΎ��?�����}��տ�tí��,-��vΎ����dl�T�w�1���C9�n�R���`���+$gv��ѥuW��Ɣ�������0V��g�â%�>=F�tF&���u�4��a�OI�q烡�+ŵ�����Z�&���Ut�_m/��h�-R��g�L������Kp�� ��MD�FJ0��8�,)�/(���3�`.i�'{F�R�ӀYl3\��i&G�WO����g�P.U'��0ܰ!�ɯڭ���q�8�5��1#f��i+%@Y="$FY�@m����e85qY��3Z�r�=��\�
T��2W��Z�O������n��ܯ�
~PT��=��L^�����)���V�`+a(l�A���ޓ�3y6�C�)�<��a_߳�X0��o��rF�����=!dU+�.����E�eHu��W��	��h��_o��S��n���r�X�;;���Yl�I�}��0�zm
Mѥ��K(�@�����h�M��^
ҹBW�:���𛊖c�MI�$K�䜶����9,���r�*x��.���z/4w�emʏ�|P�,����4�
��9��ǎ��A~��g����r�3\��k3�yT��������W�,e3	(��CI���pQ�=׮�jB�v |\Ed:u-U�ʥ��$���W#�\'��r��q�