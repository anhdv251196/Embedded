XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���%8w��X��9����C�vF������@,(2C;)��K!}����d֠���d���?]����t���5�/c�_���S;�LQ!���G|�����7������-�8lX�]��e������~Z�H-������_����������MV��gE��rᩛ�
��Y�r�pL��#Dum�bx@��ܔ�,c����Hq�9�1�mbx�8���&���0�K��g�e�@��2w8@���-�g#�'##fV��[>$�����N��I]S���(K[g����-��e@Em�D"��/�8b�$�Y�@BHJ@����Ө��A��()�jRA���h_h��Q�����TiOmƪf���~&����E��@���*���h~6&ㅠ,�@B����h;H�|�@3����9rB1v�ބ�T�}��|���Zw$�56}���X ��=�֖
΅B� ������l�R�;5[��o����x�N��sSzc�r/Ӊ�i���0��jҟ�C������B������f�Α�YN���1�q�U�i1]^׽���XN������dۚ6J�e��GW�wt;��0�֞D;�1���԰�N����n4�����ͥ��6�,�Ob�>��JA���3��OR����h�f�&B�s�z��V%[EP�>P�
�#'v�`�)N�
���3}�i���h�	���{���iA��V��đ$���t�8�����9��'�x�x�I�XlxVHYEB    1577     5a0~2��+��׀���Lɽ�1|�
��t��rk$����cM�����`m�&1�$5���u�c�Oz��e����=GA��r�#_�u�$(�H)���إ�9�<I'�/��z���;��I�m�����cRBL��?�ҝ�"EN/��-��맵���ͻU���ը������c��R�)�W.�.��	X�R{d�}s�B�������ۍ
��"���/:��Q���D+�?�J!~�Zg�1�m�+���ZE3�;��ȈYƭџ�E8��u���W	�쥎k\��K9tV�}�`�R�镲��)MO������>_����ǝ�[�'�����Ʋ��ǌ�P�#�+'�,#I��$ƃ�`�\��sɁe͖�7�R[I����� ��*�D$ݭ�I�e��3�jU���;��O�K�!~�?i�}����l�!��d?��P�&��->,���\ؖ쥗:E�>�-BL�b	����Ѡ) ���1�	V���E�.횉�&'���cm�i��;G��SnpHz�q�_����o~�Op���i
�� ���	�L�&	�c�j�O��� �����y!�a�'r�h�
�W�>˚'#��5�"�҉�7T�}���v�!�@�?��LkTe��h�2������v\a�"#�}�2���slt
�Fcsh9i�V(�w��<*e��]"~H'���CT��*��k+>�O��bS�,3��)�.�x?s�ܾ�I�Xf�m㘴��X�<�����]���t�AъW
ύ��kz�����UR1h���.��eOo@��S]�����]�3ܛA u;ǈ������aŚߔ "�m@�&����O��"�w�LZ�ap����f,���M�<9����
X^Gp�����y�̹ºaO�ά����ij�!j��%G�Q��an#��DKG���x#d9m�x��pV�=��`�@_t�;F���F����|�Y��D*�&xV>������=5��U��ۥT��A�c��k�39ߢ��eR(����!�8�7'uOSt�U��A-@�H+X�Nְ���c�h�{�\�#��S��r����B^��)Q!�q%m�	�P�m���sc�-�2Vp{}����aG��_	:���c�eE��3��0���C��uP��4��]`v0���}�ٰt���0�#�1��u���ΐ��-�~m?�l�����,c��v�Tv+��pUZ�yZf���'e�~��I�=!���ب�!A��n�,}X�<�ZH���H�JӀ$�f� '����F��b�vf��N�z�3b��y���qO=Z�C�bo���@g����ށ�H�b�@�(&�
1NẆ��|l��ָz� ��E�cT:��z	T�B�`�PT��9}�}O=?�Z�+����1���	K�