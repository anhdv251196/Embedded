XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��G�7�s¬��X7pf�&����%Ӝg2��~������=L2lO0��w
F��s1�nAe.���t¸����m������F'�*q�Qiuʡ{N	ϣTQ�É�� �~�/f/8f�#Ϡ%�v����Usf:���1�I�p�/M�������A�)oRH����Hw��u�X'3%�����>�kf/�}Q/V��.�kuV���E-~>qF��|L�,�hw��~z|j5��1���}��y}׺��{��t�[��8'��DOx�e@S����ŗe��&��aq�I-$�(xD�V�����X�+n�k�sZvH���Ee�o���FgL�~VI�^���21���H=E�9t�
c��Q�|)t���/ղt|�ۀ���]w�(^.��޿������1�&}
٦2� A���<�ak�6i��r�c�j"���q��vW=F�34w�C��4{K�C�}{#�h$7�%�urA2���6K����.�����S��E�S�8���fS||ǡD�+�S�'�D�/$]<�+�|�U�����4/��o�3������dg��ϸB鯱³���^]�����o|gH�����(1l;����X�~3��|����ܣ]Ta�D8�J ��(u��rDN��EH�8G)�j�AU�H�? �x�G�g��M��BR8|P-e&%nٽe�(�^�/R�V7�=[ n*�a��)����Ƙ-����AH�?YV��Wv!���ɫ����R��t����"�������۩XlxVHYEB    1d51     7b0z�:5���rv4�>��q�0qr�I8�Ȳ�j�	��s�ZIǍ=r�<w�x`��P�C�%1��j!�]b7(���Ar���Jt�o�5љ^R��>�)6 �w*���y��e����uF��PȺ��h+���ɸ��v��0S
��7�?���,�U��
�	��r2����T7�*R�sI/�-��:��t�czZX%��A��/���|������]A@ s~��%�n���e��T��b_�H���q����?�pB�ٶ��k����&>��L3RHDQ������;M�̊�Ͷm�e��GKq�̢����Ψ,z�nG�HM�ǘ��#t�-U�d���H ��s������5��^xljNvyR�i�0�,G��:4M:�2�/1/}鹷�c�zSLlb��L��my�۴ �+/sp��N�k{܅?�a:XP�h.�H|ӳy�р�p�Xof�@��|#LPbJ�H5����R��)���&�}�%��v��Q �����1�uJ`f;qUN��. l��@�t���Xv�ٟ�s<b���ӟi���o�I#�����a�E��c%�&_3�@:Φb�4ͦ��>(�T�C���	�*`[R�����v������ *�=�M���e���(^�(W[�G�(���lf���� l�G��?�Y��k%q�.ДY^)g~�J��G��������MT�D��\�	b%o�q��8
w�ao��H�*=|5�b]W�zp�o�eO;OWu�[C���wE]��r�)�Թ�A����b�A�~Y�7�b��.#F@��|�hc�[ʐN	р�Z��tJ��2O�b��M�0������2��O,pX�#��B�Al��c�k�Kҵ��x�6Ay��R��D�!�.�ǐ�V���O���,���0�B)�I�9�hI4��������[�/����rg����|a�������ݖ��^1�駜>�L��6CT���x��@Hi�R�nCFړɺZ��B|�U�5��׿Y�hl�=�u	��fn�*�t?��5�|8�j��rr"��cw�	�k��*�5�a������1�%5f,��l1�p�����P,�.>__�O�0 p� ��ގ>�����]K��µ�`� հo�)a�Ą���R��uU-�H y����
��j1d�"�%��W����w���rHh�r+w�:�d�lhn0�t�W�w쿃*e���J�Bۅ���
y	�t��C��⿩|��w��ڀ�XQ�5�*Ɉ���͒�JN���S��t��wkk��wnb�i��Շ�m~�rn�L��[T�$�{{P�Y�	/9�ulQk��F�����; ُ��>�aA��X+����0e_A0{���5$��a�������6�B$-�XƋ0�����W���Ԃs�sT���rĆRZ�����(ʝS`��LtF���0��R�d1��<�I�ݺ|̅�߽������]%a��Y�Ҡ,�ʘ����Đ�h%�xW���}JP^��&�1ꝥ���%�q�;=�E:Oj��M'�P)�3�*x��͒���ػ�i���(�t`Z����d�v�(B����e��=�F�8�;\�=����� v9
z����/'�(�B�%�FLK���^�]�c5�3[�[ԫsz^L4����`��s��Q��0� ��A��f������XZRA��>4E���X*ڴ��]�YY���L�\捠.���&&8���C��L�I�Ǟd�2�-��Q
��V+t�{�������Do_� T�_�Ѐ$3~��vx�`5����%�7k��߳p)E�٘�����-3q�����~zW�롛��
OV�!L�b����S�k���Ur��IIÎ ��`��+m�m��}@0�7�� E����'�%�bB���-U��餩��hE	���տ����_�M4ddt