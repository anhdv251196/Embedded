XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����]Chm�$܇A�:�,�L]�/~�xI��A
!vi�p�Lbe�D6�[p���`�:ԝ�ps��M���bF�Ś \�H�g�!hKT�>�ִv���BC�aMڽ6�&럞��z��·�9�t��"�J���9���B4sJ�ҁ~��k���du�����Q��L�/E0��i,� ��T����`v!:�tQ6)����-�yŢu��O2��QH�~c��a�G�I�V��dӯ�i�Jx�L�'mO:�~�Vv_b�H�Q~�������䱻]=ȭ����fT��$�ߞ���GM���w�x�[a����������B��$���
|�)���(NAd��S#RG<|�Q��.�A���)lP\��ԇn�(v�!�W��ߢG��7�NQ�N�^Qȱҋ"�0���R���'��t4���Η��������w	�R�����߉�a�
�/��"���Xa[�ܕ�`�B��j����v��8�g��Ȕ0n��l�g`3ܞ�\/#�i/��p��Z	��p�:��LQ�D�9l(�ԅ$t�a}��KA(�BG�KǮ~
��H܂yӰ�Z"�iE�FNh�BDx�Ǡ�$p���<Q�K ��9�`��8:���+m�Ue��X��P���(���Z�Dn�*������ �ΔHp���U�Gޔ9��gUVs���e�|��@n���^�)�JN��w��wZh6��J%�r���$8��ԛ�o�$�잒wm9q��F�����XlxVHYEB    1041     4a0���P�X<Ң���<�#�ф	�_��E����N���⿢�%a���=��9s���G�4�q���7i�y�;;��|ug��m��[��GД `�$���E~a���UP��#A<�<\£���R0SXm�����Ȋ�x�\b�I����
���|6D���]�`�u�D�7�sMc�2����>G��J�^�թ:Q �!��a�3p�/g0JZ>�����Go���b�ʺދ=v��0Tzg�eB��#�\�G�n0J$T�Kd��!�4������@��,�a�"�R�W��P�h����K���� �c��N�A8!tP��l�\�:HU�>�q=�ݛ���S"�6 R������"�6�6�N��y-��,YJ��b�͕;�4E~�П�z���l��!�+���}T���{�hX�F���G/T��]\�7��3j�M�ʢNU<�N�"ܨ�a�j�)�X��xf��}�(��0�4� cuxs�yFA���,%�6�a�Ǽ����6��T�ʣ]X-E��w����X�ÿ��K�F��W�ڔUqլ���O�$�Y3���Tz��t�ܼ���W���z �k�Z�V�KN�	B��g��`���/�N�Y���L\��2x<mS�N|�yF���C� ��TQj�v��A�&����!�ݒ|�lg6�s�Z4`��}ڋ,�����zex�Od������P�E>���\1���2�ޙ0�<�����.������.r�q���+�AǦ��5�`��N�䁂2Gk<���Պj����2iݬ���ig���pWr>��$H����עq&�l���Ao<;��������Q}V����桯��V]�#�X�DFV�}]��襕z����Gi��,�e~W���p�]$�.�p�#�M��}gfUT~����=��H�f`���D%][t������������Ud�����Z�T�KRY��z8FQ,���	:{-$܍F�{e�ҩ1XT�w?Ѿ+Z�f
��e��)����ԯU"����-Rw���	;��������g�9dFNMda��E{�+�K�*�]��e/����#����.��S{9�l�7��Ǟ��׈c�"<7��+\�#ɇ+��/�P�� K2����߰

aE�����