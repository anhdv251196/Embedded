XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����G����lb����g���sq�$تh5�|p ��K����K����"���q�v���7���7�Pt��5��@�Ub[�IK���*��˙6d��e�N�%�R"u�8��Lc�������wÐ�5����d
Ԩ����C�(��;�O��Á�������ϝ&�V��f��/���Lme�V4�2�k��K=J���������8�,qT1��[|:�qJ&a��p	�y�o��!?� �G���p*�;/�w���$�nl����{����¨����1�!i���m�~�O�͵A8�>�\AOX%�q���>�|���T/Y�������7&��D8#����LIS�<�(=ϵ�+�H5䮩!<yu�c�!AJ���
�O6��+3�ɦ��	|�w_�q��ڐ����R� ���F��f,�~�%|�����4ո����-wP�x��o�����V<N	�X���^��=	�J*+һ�7��ۆ����űnűG�@ }�"��+t�y��n��*sg�e��P���ʦ=A��tÁ.� ��:*k
�j���Y s�'�gwA�w���G���U�N����(���5w��x�2HoW��Ǿ��P�kS9 ���g��W�|ܭtC`:WE�JA��8����-Ψ��i� 2cζQs6j~_aj�#%���xxjD�Z����1?�>)$��޳W�	mCѩ}ƣ�/���>-���� �n��K$L8��1���k0XlxVHYEB    4a09     920�Uxʤ��Y/��'�Kc�LB�QX`�&��_$b�aVk��w��M�kB8�����I��4�V�.pB���+t<���ݕ'�C���0sֵ�s��z��1sQH`�A��
$����ӄVM��Z�È��r��yd
Վ��A�㋵c��mV� 7��O�����i�㡖Ŭ��ù�
�ǎ��/#T�/�[bq1����3�� �:\U���+�gO(S���B�v����dq�̮y��@��(�$N;d��(nQ�h�b���ԭέu���Y5�!��Ѓ\�,g�1����[_]9 �a��z����^��T��E���������9���ro���x_>}z�]/���?qZ����5,6M2���Y�����
B�����X[L��`EZɰ��꠴��Ot<�C�-a_8؆G�:1�]=�5�*�����,
-���_��-zǵMڝ;�X�>���K��.��Z��(���&\\�{�%c7�7��Ҕ���g�ѣm�/>���c�r�#������*
x�U'\��랆�y�q��I�������^�7��Usƈ�����D]����v�����?��Ii �_��<D,/^d|���d��Ν���t�	i�j����4�U�8f�F��q�a��<�bd�Mڲ��@ z!��"���jط���N�Ȧ��[ �%�R�A��¯p!�A��� H���>��q�:�@������`������Ͼ�uF8�=���x��]m:ͽ��Bh8XL!5�dP�8í�j	��Y�Za�n�|�y_�	4-��8e�c��į}QX�9����g7��i�j)�V3�q��'�%@e1ZH�=�&����T4v��L�Q�_5�˹��@�M�2�7����	����Va�)�;�b��uBR�`��d���X��1	�-�~M�J�G��>�KM��� "�3+�ؽ��w����5IN@ ����冴{D.�w��#rIi �	�n����af�l�hU�B�$(%�`�{<��[@8��!�#�9�{�ۢb�&9���4ǐ7�[�Dͣ���<���%K
Y�-5��F�����[�����X4�B�/��C~L@��o�y\���c�=��� �]������í�b�z��0ؔ��1[�r�y�SyA�N��d����*ő�T�'Z���175��h��Q���͆�"�lb�Tm3=�\"8ÿ��"^��b�C@����aIE�N!�z�߯-��o��H\����\͓>�G�܈~����2G�?b�z��(�2����)�����(�ޥ�Rh����H~Ub>��-�oy^�3]�Ǥ�?*P�#���
����Q���t���>`H�&d�kl ��(]�D��^9�	q�u��Y�d�5"o���m���b�]�2�mw�|�����2�Gl�YA�w��xV�j���#}D<�n�z:Zs~�}Y��^.���[�����e�h�L�i�\pd<�%��\�g`���W�Q�7�s*Wm����Un�$*-���˵��c��f�e͈�D6���4,���{���y�6FΖh������C��Ӳ�٪��Bz����JU+<8���p]+5��Q�1�gv��IēP��)50��X�d_�F	B��R-��T�"l �� g�Q�u�^��P�G<蓊[��[�>{zK��_-�R!�&��^a�4� ��a����U�o9�ŒI������3��A�Ñ*qs��RH�Z)T�Q~�ڿP��hNm��z�]��{z5k���f�f�v�I�~r^vE�� #G�֘�$�Y�M��Lyً繠h$�k��ޗ��rWg��v�u�rs�4c2Q(AlbMv,�`ݐ��F����4�D1����Ɏص�w�9ȁ/an֝qa�[-ȴ��G���<q�-��}_��]��u�yxI�r���uA!n
[�H�%���]����\���������1'��o{t(�*����$ϡ����~����R7f��K�A�d����A�C�鴌���O8D޽��g���Y����,�a�E��uD�Ur�:<�<r}�����k�g<��v�~Z�����&۳m6w�'VI3�	�64zr�ͳ����&�i��v0S�>�͋G��0�&F���N<%�X��u�(������C
&��Dk��ç�m�lIx�rxFa;'+�	�n�Q�uD�t��*�f�U�l.�Ɇ���\�6�P+�X=��~��0,촙���AHi�=�/�u���םlMA����#�[�1�7��И'F���ĭ����QJ���^-�