XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��������~޳������#�YH6��2�z6��G\�>X��F�����l+]ߞS�UX���-������H�h �ٴ�����Ҋ&�zYX�b�B����s-bŁ�g@��M6�e��=uB��-}�m���I�^O!����_/�qSZqr�]n/�ohʇΓ�m@�mR�Q>--K�8B��;2mp>�Y7��!�!�N���7����V�׶v��Z�n"������	7�b�Wl% tWj)5|��{�>Bq��q��FT3
���A�!�^Ű���PxR�mlCF��۸���H��2���j��8��#�`��X��옱�O�����Ԉ�ؚ6�#�$&feq����g��A�;wDXܘ���_i���6�>ḑ@S���C���xR��yA�P����j��|������s�$]ܼb��W�l�Z�_*��$�N�P��w�$ I���SRf����@#q:}�MRT�,Z;�d���3Q�r�E�iZu�}M���ґ�V�2���W!�s����ѣ�!�.�Pz�b���b�ϯ���tBqr	���/!hEC
gV`:���_"��b�\B?J !����n\�~'��f��0��a��7�0��+���AB���WĪ=��ŷ��j�lZ�X�ږ:��ٌ�<g�: Qo��6��:��ȯ��-��'����A@u��8K+��fa�寔^d��2�ƭM K�:R����vYm�*;6�F=X�j��O�%��*-XlxVHYEB    9b67     f50|�N&5z_[��N�뼻Wc"XOC�4�������Bu���?� I�w�J�5u�	��co�|b3R9�-�yB<��*����r��N���X��i�V 7���\"���51S2�Hc�4މq��OT�yϓ`�"�ȹ{��;�
�N�[�Ss;���dF���э�4J.�<�P��Wq���?f�Ʈ�&�2^��f�2w�O#����i��A��q$i�u3V-�0��2>���S��3Y)��b�m.��0_"?'��a&���ČU
��〔"�J>ߑeR�(���j;a"�pG��;���.� ��ֽ������������9	^-�TQ
�	{2�v�ar\�]�Oc#n"r�𔄵�w�̹���5��!�F�1t]�l���]��u(���Q�>ޣ�y�~�)9��?p[�r�����K�����*C��	�xߜ(7ZƊ�k�)���������g�%hVzl`���#7�� $����������%��;($�o����W�0�_�d��6ڌ�3)�����%ƇX��
���X�����w[^; o�u;���O��ۮ^��u����$����ց��J�?�� {��k��-�;U����Om����1<��:���C^��ᝄI��`��"Z�� �U@�uv����P��E��f�)�7�2���t�8�or�P��K\ܵw��f��#{;z���`R^����-,�����#�Z�D^�(���D�p�*̌&�o�5*6E��,�-{��2�bA`7L�~H��m�p�R D��$�p>�&�h�D[g��a$>�[;b6��&������
��#t�$菴��܂ůG�� c���&�qh	�Y�0pU�=5(�ҹ��0�J�A�S�v�F��P� K�	TJ�&�����or��h��_�i��p���m/J��f3���s{��4+��6:��Xu�RҒ(ç��tAGJF9�N�{�X�ө��������}���f吖�z�U�H��bxi� �7phA�G
So�W������l�|P�"���]�v��5�EM�o�$��t�=�`���@�m����:�)�(Z�G2���Q�p� �=6.�ɟ�~!<L�����*��p(��
����G�@���_Y�P���_���v�ؿ���]Q}�4auZ�s�9\W�]s��ר\
�]��xTv����sg�V@0���{΀^�H��;�		�*��S�8{l������*U�=�}�cV�"�Q4�i�>Ď�y7�y�L��n����*�f1��N�P/���H=U��zoJ �����ӻ�]:�\
�o\�]���P�"ȇ�z&k=�#T`&���?tX+�U��8��-`~X�n���M�`pk���p���UB�E+��-�M5�����(��6زȶm$�s�-�~Ӡl�F�_�97&f�ܡ�FO��寿 *n����%�� M��]J��cm�^�����]�.7�Փr��'�8�r��(�=I��F�Xw�L����$3�U�U��'D:ᬭ����h�h2Vsx�ÝRx���Q�ML,�k^L�ol�!�L�E�ݴu�2q���#5/�]�!`�
��`R���u�-�ߟ��A��%i��4uP������̄0X�39�X�h��1�>ؘ���;������:�.B0:rlX���+V
���嘐re?~ڝg��2�����Y��+������o���,�'�AZ���aӎ�G������6���~u��P�pMn��jRꮢy��u���(-n���F-�G�+�Ͻ�΃��,��^&�*��<��,Ŷ��������ܐ�(��7�jk�ť����猔��9=3���<���7['�V`��%Hi�p�4p>�S|8�WU�C[�V[��U��i�.#Ot@>/����7K�ῷ	�|�˝��XhC��7��$J�}{ɒ�aF$�nR�"b�B �"�`���]����Lj��Q����R�'-�����1�jC=�>!�f���2'��f72K�eD��̂�FO���h�.�&Ec��@n�k�QEp���D~�w�;T<�k 7j=��Qx}5%��<�5�'�\�r��V&HI�N/���q��>y��4��SJ�W��<ܦY�xZ٬*19r����K�$��6\����q��b�4$!Lr!���n�pj
��Mmՙ��5���v�e]T��=�����Ĳ� ��\�9�pv�����~��R{⼆!�#5>�5?e\6����Vx ,�����<���<��t�֎D~(���űJ�����@'cK��8��X�C�������O���G]W��\��7���ړkx,Q��Vg^��\ʰ������N�,���+c�x/�ց�c�'%��W�g�%֕݅�+Vҥ�TBò���i�'�(��NA�u)�>��p1��#p�D��2�F�?t��3HY�з�(vP��c�QDi���Hv;?P�r����GD4�֕a*}��3������y:]�2a~�)K1�T#�N�"�P��Cc<zrT �d�E��(ե��6�$�����#ª��I����sZ�!4+Q�=U�BW
`�dﱬ�E`��p��Gv�o�w�Y1�q�
�O�͌�n4j\tF�@����v�ژ��W}[��U�q|Ϟ�I@�±u<�$}	\>��:� �&��b��tx(�)�2Dj~f�Z#��Б�;����6B	�U6����X=�~��@���o�����ܬ��c"�t�F-H"�Hf��K���a#k'80�3
�����aa�.�J�'�`�?AM�UK���H�-�<f��YM���o�z�ߺZ����2���[x�E^�6˫�E���Nd�p&ab�����P���Еs���%Iy������l��G��iu�� ��<�FG�!�O
�8p������M;��%�P�)?�؞܈`@�a
�|��q�Y�%�ͣ��Բ��?��Bk �g�V��.�u��@��t�J�B��YC���`u3=i6�@B��uTCڊ��?O{�yJ�2��<.�ﱸ�=1��gvx"�}R�]�y��}	� FiVW��I��F����'$�~> %1��~k�П�O�<�'��
�����/ j��FB뫓
�Ns�H�e����lf�V� �a�w�A�cޏ��W(Ϭ�+ҞW�=��Y
lc����3v����؉9[)nuunnHB�l9��凲�O�k𗶵�g��{�_��v�Y#)*�L�;�F��iz�Y�]�> 4Qp��w1�7�^�k�ޠ��Ƅ�У{9�4�X����IvS�ۥ�S��]���	d�����SBvm��T�(��o~΁�|�n��>�g�"P��xcW�a��/񉕧�3O� �w}쟤K��F`zmq��L ����"�2f5 �G%�������Y~c�J�
-�*D�/��@��	��ų2��
kz;�dǖ������@��j��� ���8���bK�~�l$�=Ӵ�}#���q��hɀ��ޑ����T3��d��E�N\b�bB�7��x'^�1�B<�50?�O;{PBK��&~�q�����i[�7������� 期�s�Y�?��	z�vbI@iL�${������W��`���O��/��=�#\B�X�b7�߯<m�G�&j`.gk�a������H��
T�{!��d��K c3&��fa1�O��GDH9�@�n�>w�Q� �Gś�h�펥(����$V�`�T�d�oz�w�ӄ�����m9��V�!��|��8-�f���b�O�D���,��D¨8&��2'5U�ץ!�I\��f�N�;5J�ԭ�v���.�2�p]���"͢�w�]t