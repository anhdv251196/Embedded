XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���OHK�P�(`"��}�l/��8��cGJ��,RQߝ�T��R�L�8*���H�	gbir�w�oj��U�=��zE�����#$զ�}OHW�m�3�"B�8��V��7����U�r�s���o���L<�0�:~���v,Y���*��4�X���h�J�jv,B���݅����3�l�������ԫx��J~ C�y���VB��h��Z>�h�e7���r`�0�l��f�+��{��Z���EF�_�f��6b�mS�@�KxP��r�YΚ2�s̟�,�`b�����뵎?A('N5�������Jq��Lm����ʨi���ni8��Û�!\/�����nQ�z�f�
 L����l@Y������f�F�#*��*�P۬۠�ɦ�N���RZ� ���f�~��	fd�`X�wAã��JH�z�l	
�1�Q�� ��?��Y���t�EI�'�c�1����ެ��#괂Xh�w��{`�;?+�i��0����o��D/;=�ʄ�n����ԍ��ni�F·Aě�!t_�׹9�voҁ=67�-�86��/��h9�!Q����`}8tt�n�.���ca��BԑQv�)R���Vb��Cz_E5
{��MQ2���>�V�Z�G��j+j���M�z�FS�'�h��=��������֥�0o^���M=�߄T��6Q��̆y�ۺc-p�o~[�r�H��b#�b�G�����U+��m�H�r��.�������FaXlxVHYEB    1047     4a0���%��K<��r9���z��6 >�Wp�\/��J�T俳$$����+������q�_��K˾�ĺq���'��[�U^��e���w���5XCe}��c!�{:��7��Ү+�N'�;��=S���8~K�<��X����0k���V}�,�K{̖q�hy�s��C*y�U>W8����Y~ς�wf	Ւ��]
U�x+{>�^�ox4�=��'�Y~���� �ߪS:Ȁ��̜,p�<��I���C$��٥R�~�`��G�(��w�с��c��_�XA��Ai��!���5���ࡃ,h�9��-�����~�.klѻל��!��5�U��UN��I9^�%'�{D���R��ˑ��iZ��ru���`2k��g��vt��$[O6I����a7?�BԮ���*Cm.��4i`'WA������m�[�ㆬ�`c���x��k%�c�t~�@�Q�^�G��^v�������~0�
��*�z�J�z������WQ�� J�h?p;��OPT�A��E�1P��Ņ�T8����W)��<X��=ӌ�a��M~FK֬����o��5���R���C�>�8�-ʌ\�s��X&���qX�'Q��s�(����;��JmD
3�`��z�^U]�6�v�c�9-[���E�c�at�0���V�K��*��C���!����o�0)��Ȃ�����N{�Ǥ�*?G%�b�{*y��K`M�F*���l�sre����Q�HM!-��j��PG��z�2K��ݥI�0ֱ-c�;`�IGE8��z����%���E��P	�J�����k��Uk�1��G�~w�s/�	��=<� ^�0�����mx��p�Z3��[��-��ET;����?ܾ�ӒN�Q��$y���a4߈���k�S�����E�9�$���(���3+Au����f�m&��.$���?��o�1�%s�@W�_V0���-�SߓN��J��å��}� ����cz�T�ZV8נ+��86��$⛞|!��q����@U��*�}T.+�g�d����)�iDWv�t�'m��~�1lu{����HAd[+%%G[H�0�׍,|�^{�ѣj��cs����N��G������$�Lj[8߄+>�2Äu�yaQ�	��娌I��H{}��%�J�