XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��;�괛�hr�-}*���r��2��7A,�]gWuK`KAo�,B�"������1~���x@��1i@������z0�>��زŷ���,��j�r�ߔ��~
&e)�B�ޗ^��,	��⒰�4�4���p�2��^]���6�9OX{G�?ڹM���c�5�jlu58+x�m�5��n�&�R��׹�
] OO��{���n��Nv1���"�aD�(��B��ddi��v�c�@�����;m�f���̏���uQ�l��۬���3P�#�QȲ�)��8ap+��Û�[m��N� �<���7��h�t�C`���q����l��|����h��@q*HS��ڡ��M�Z���y����GF�a�b�A�˨��*�y��9�ӽY�oadx�I��8lp��5�|U�2�L��Iר&��P�C6���M%��L��P����?��؍l�H�K/�6����ȹHC9��$��U�H����c��	wP��ʡ�Ϝ�B������M�QwE�ZJ �ƞD����Q��X/��8fW�A5��i��?�-��P���4I_������p��YGic,Ү��!��7l}@�ll�иOu�3�He=ϣo0%�/]R�N��#q	�}��f���>�%@9L�3���R8^9��䡴�}`G�Mޏ"E�O�o�L��� �R�a�v��t>8���(3y��Z)g�@���2�Rl���pS�T{�3 �fZ���ɣ #�*M�[sa��`=�o���P΀��A��Px�J��]ՠpXlxVHYEB    1b22     760Hh��w��f�J-"c�M���	#��ܸ+&�c&��bR�������!E��h��?V�Jn}�ŏ�ֱV��:� ����HRd��ɬR��p�&�]�^���\�����V��$ϡI��;�����j�)�k���`��oٷzOz<A@�_b�s�l�ϐ'���`y��/�m�b%��5�P#ցoI��w�_��b�3\X�;y���e��ͩp;z�c�M�U}9p���G	xƞuM���k����U��fw���RH��>	�{�S��rN���F�U�؈��q�x5o�޼9J��|g�Dez��&|�[J�~������������6<t�p�"���Hǐ��4"��+R���[6S�h-�	�֬6GC��������7���=Yv��:��D��Ri�&jn�'�<�g�Ot��bii����Ti���\&��}��/+׮��|@��~|�ʊ���w�7sy� ��+;�N1ϐ{���{�p��W�F�w�L�Ӫ�C��G�"��h�+b[2ra��L�9�ܾP�s�΋��߬k�o;c(p�����?.V2�.t�M�����\ V$��-r���$�����v���V��Hv�B����b������@��h���.z��fS������%>_�x�t��<%[�r���&�
F~�`Yw�+��ݹ��#�U0�@7ww�vz�U<��*�	h�4��=��<<N�5��c"e�]�p���80��Y������\�6�~��I�Ā�Cv�� m�nP�tV��r���߷�:��������6(��K-?�^�e��i\�U�
%�;R���c���g-��E��UY-?�)s}�ҍ�jT�'�����Q=���<����$G�Y'�YRk`�`��-�5��4[{7+D���yre	�|��Kʥ8���Ձ�2�Ғ���s�O]��9���5Q}��5�˄�=l�Mle^�g�`�|�:Qp6^b�cx�u�3�G�0���6`!��#B� �|�e[T��⣫v`�'��-X*0a�a<զa�93�n
%W�����!�Bf��;����\��E=�M��� ֓	���;C-0K}�+�bs�AC�M����"���j.C{�ώ,qm�`ީ��K��hWH��&�M�%�L�Lc�Љ�/5����{Qy��#Ȋ�$�����O6V���ȡS�&���?|1YF�L/�_
C��4�k:kcI�m��S9���G�[|�����e`EO\Ի��$x���||�@ c��?�v�NF�^������%7�!�ܲ�f۷�\y��'+T��j�)��Z]4��RC�ٱo����-�Z�$�,���$!��Qj����M�,B�y�b�q��i��*��c�˨��#�5�o�A`������1��ڪ���x�i0H�r�y'n�'�9�d��M��tj	��)�.��aٶ9X�=�V�O�zJ�!�!���G-���NJ�6y�Nc�X�CCJu�|w��,j��V9A�ZP�VJ�ekl���aT��N&�±�+U��ě&BO�۬�$��"`��F4��L�N��7�#�T��u=~|�X�f���N�9�/섷*'�{0��u�b�u+�q�i�loKX�t�~R��)<�te9	�?�{Ȳ��$ƽV���W�4I@�ZF�@���}NM*�1#-��xl��t�����ۧ���6��(u%�U����"������й�^:�c}��P�oK��[��A��uÀ�iI������g����[���;�J�)T�����<q��ZlG<�U���rZ���B�LU�l��;V�}�)?W
��*����J�>��"�����,l��*�l��4���vEY