XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����[C���>��!����̤F&_Z6��<���#qO*;��l-�n�F�PiE�J�'�2-<鑙ؕ{�8�������3�s�����#�;���XC�F��������J�+��� Ɔj�6�o@ʶ�p"B�����^�;� �_���-Fb�B�u)}�.����"��_Hg�[S��d�ZY��d�Kl���a'�$�4b�-�(G�������$�U�Ϊ��Mɦp�ėNcQP ��,���o}e5�"=y'��H�v3'�<��f�I)cL�r�=���H��AT?�� >d��I���������&g�"I���n�I��x&h.y��w���ѧΟ�uPx���O����Ǿۜ��/闀�K:��yr6��Sg�M奊�j��j,x�0�y~����lCfL��a�H����Tb팪��[�����Y�6��,�酄��o-�h\�J�@�� �������@O-8������5Ǻ��i\,�*���u/�_!߽Ot!��[	��v������*���z�޷�
(ļ��=�`��V�͉�Ȧ�}(j��1�L���C)]͝�6�Lfזo��v�"c:�q�/X����b��N>����qE�����Y�n�^\6BK�/cl��ާ��9�$�654ЙuY�y_!������	Ǖ<BN����������X���' ��kM�Z*#�h/�[>�!�m3� �,Le����Ph�N?@CG/�mȻ��Hn9b�'JwXlxVHYEB     748     310�B-Js^���o��~�2��#sKԈd��EвT���ȅ�P`j{V^:��iRpU���c��;�3�i�.�{5�H����ɒ��o[�N�$�yjջ{�j,;�v�Э�6�o��Ⱥ	']����ᬥk	U�,p�[=/�fz36��w����T�w���鐂����Aw O59�E_/�gƭDt�=��V�a2�VϽ���\�H��( \�`,��D%�w�+��غp��p1 }�����o�H��,��HQjo���L�pP���z	��7I@����<[� �JVw��8�fU�$��� H�^��#v�NK��$�	JF4?6e�0���1G��ICQ��P��S@�t-F�w���?׮�
���|���|��<OA�pxUYO�&���2�v�S+P�9��ϩ�@3p���f��mz�ߕ%�vD5$��@?yA/:u��� ���A莍hL�1p�K�Sa�T�b��%ζ*e�%�́��)R-x+�d�>_wL���E�T��rQ������]�տ�{��x�͛e�3��Ow|M���UlnT:�4U;��������_k��i���y�K��h��[g}>^h�ծk�j� �ɛTi؃=*���^v�~��|�^X������~>�c�~����I�ܷ�=�	�-T����qQy͊��?S�� �� ���i܎����Îu:��S��z����GTLn|�W%e��v-ڃ^��`/wQ,^
ɂ8���B��_����zrd�HENR�