XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����1{��̎2�q^t�^9 '�C�Tl�m/$�x�z��'��N������H�@�����X�:��GX'[�eD��>ގ��`�O���Le���]�V(Z�.��!!���D7�M�tJ{<ĊV���s�2��&��Fj��h-Q��W��xЈ�Jܤ|���s������Be��|��o��X�%8�O�ߓ�\��¬dP��.$�@�pJ3���JM\�@1� �W�4[���n�=��t!�l	@JB�ۗ�
5�1�	���q�����e��ɖ�n<R��C����|�&�*$L��9K�cף�*��G�h�q�DhLj�`��?nab�z�ۥ�`�4햹����^W7���a�e!t�)�X-�⫿Q[�öF�n	�j��2(M�CO�:��N�3��퇛<�V���������v>>'�G)��D�LD�(��:�'�@q�|�//<<<��6�M�@�{<ک�~?�\�"S��+��5�"ҁ���q�C�f��kp���I�Y<����G�~�~I�Ϊ�?
���G�v)�����jj�~DY/�O�����:V|��:D"-mBVd[��C- �������'
�z���+�6�������h�Ĕ+��Č�7�d�Jvq�6V�T1.��G�^S�[��s���.��R�~p�iX�AҺ�i����< �{�B�ƪ�����v��˾;�뀄o<� �Vےj�䋫G�;̇{��e��a�#X��2�����˃�	46�AXlxVHYEB    3a1b     d40��ѽ�yZq�p�!�̃k���\W
�d�!
:����>"�e�"#�Z�=�A�Q :���p��x]A(�R��C�4V�Y����͒7�Aʪ���x�2�Z�KZ㞟��6�p�� ��R��+�����ò��R�5��T�j�9ט�6�=Vs�:�bd~����I��j*r�zS�:ᘗ½����o���D��c4�db*t��By�4�Ӏ����kj��U���	�CǱ!fw(/��䒛�hZ��n����0����㾒�T��{��Dp�:�ɷ��չ�2��9�ώ�{�',�m 0���/��$�; "F�:bͽ���B|0���f��a�5�Z)0���,�)�>�V{ì{���,�N濑�8Go�����z� ��w��
�����Ag��`I�#���#�:,Xg�Ἂ�&���!;H8i�~�J�`��,6�D�Z�n���,Ytb���1��Ep^h�� � ��<ʠ�ɍ�)D���vt������?��X����H�S#���v'��<�"��V+L�7S�㰣|���.J�jv��A	�&��/��O01BOըde��L�k��������f�4v�	;��х�!~�q�f���i�x���H�������Dz8/��U;��-�N�Xl��M��@r�P�����-�a��U�w���
}`��ۘ�Q��c!�����
4��D�$ã�K��mŽ�@���GD RzT��<v��k�j������!�-��l� � ����"��fK>��٫ F8��K��5�2W���}��P���o�QY4U-Vt3J@I��Z�Kѣ�� �~C���n���̠N�C2�B@Ӝ��Y��2qŁG��&�>I�!��範%nk|��B���z��9�U\,��Q�J��ڧX
�	��1�8ze�_'�\�M\���AY�~m�YyP-aPH�3��cu!�צ���el�z@����eF!�pPJ�y����0n�ҙ����8��/�O�B�P�Sk�g�,�����j>P�z-v�ߴ��겢�&iv��K*�A�fH���j3�sh�	�,��7yբ����! ���gI�Y�c� ����b-�H4w��<�]����H�E @Z�f�O��8�8hJ;�v�9����!OM��o5��#�a�h̠��ًs�s�f���PKݬ�2����f Zǿ����������B���K�>��1�R������z��[E�`��cx2h���J��fHNa���]�'���~%8��6���p@����vF�5�}��el�n��|a�twf^��G#��u_�4IQl�/�I��w������&@���+NiS{�ɽ�ۮ�$�4Yi[��|���M�~�P㇘�7|)=.�
f^���
xN��������_꜂��_� }Z�Z�;�"F���{(hT���d�|��hk�]��#��'j]3����S��~V�]���	��XX�>f���k H�H�����zwF=���l�a!�Ol��/�گ@)Y�������X`O���f��|�-�䨚�y��}��������4�Y�3e�6�̝ ��f�a��aV�E�-yW�����k�J'9��U��>M`c=�.�Q{�g�6�d�<��i�<�έ�\��e�J9��^���^	5~�/܂��m�T���G�*_a�~�c�
R�Q�xjT8͞=�s��֞}��D@|�F�&]�gqї�"��+�� � �:%|;q�4���?��+��:��Ro?�-�r�8�MFS/ː�E�A�;��+<f֧�Gw�x Hw�r�{2
�mMu��u�V0�&�w(����WB8�q�0Y�1����� !`�]����6��e{���Hd�lGg�d\����7��;\���L�$�#��7�տ��<���)����l+����7U��ρ�(�ѩ]���2�^o��B�ꬁ�SՖ����aW4X:C�2��A�e����b2��#8����(k�o|�MD�(�Ze'�B	�ǽ��)V�,E���������u4��U%4os|�Tyw�vjiv^�w�uM����K������Nĩ� �ݦ�Pg�����dzIS��|dF^��������w��kM��b���uD�+�(�gjn0�U� ~��\�k�H�
i�}K����H��j/��J�_ W�zn��N� u�*{*vb*}�����|���J~�G��;w̖�~u"��F]����O|�j�M^��;Kٯ��� �03��Z��n��Na]�ك�7*��Ցr��Դfؔy�^�1#z��]�E^���ī��U��`����Ce-ظ�j�@��V��V��,d�0L
|-�������Ǎ�P)�׊r�_9$�w�lq�5LE�]�_� E�jcV?߭�b�����'��m��Z��=���g$���=jK�s�S���ӆ�+�;Ȅ(�#�{��UK���s��Q2���?���/��>�q�^Ő0o��P�e���u'�u�A5�C��դ�8���=��'?g��+����q��C匜7�}'&��{Z�T���GM� �6:�1қ��R�s��*�H�Z���V�ݩ5�#��sB�E�7��?W,�<�Z��w�@�au��W���u���>#@2HU� Lf8oՀ����Ta�el���a¦ncj���m?��I���o�ͫ�F����q��)��mUl�jP����E�G���U��E�s����#����û{؝n�b�F�l9����v���¶k�������S����ـ�����G�tØxn�v���{���4O�������(���9�PY�y|Zw���1@��lNy;�j��e��e���	r��Vj�^#�3����F.�vq�M��m;)ys��jg�p�g)+oF�/O����z���1�3=r^��f�-�����i|Z���&ֵ�ޮʸ�	e�hܽ�nyA��vD����-�����5���v0W�V������p1�?�>�2�J�{|+w+}��p�{~�����ڍQ �.���x���Wx�\��^� L�)D��4��(��8'��4EX�rp��v�gwE�d<9=�#�T��Oy����[Ԕl���b��#f��sL+�(
�a��^�)�'��E������aO W�[nTp��f���*R���s�h���[3uHNa���Fx_nK��"q�@��7m_f�$O������ҁ�KZv�c���
p7������u3{Z�Oj%!,j�O�W<P��.��%h[�@闆�����JB�f��	���`���Lx��x4�u�.Us���ֶ]�m�#�,��z_h�RGjm���z����w�,