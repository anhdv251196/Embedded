XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��A�f��Տ`��h<�k�`2��R���w����L�������8 ��(�գG5	?��٩�y$�#V�����uJ��c���Ӻ��w�����;�^ZL�^ޝ��}X��X4���N%��,T{&U���moK�zn��+	��ж��T~�ǐ�����e��I��,�]�3�:z�c/����S����/��BcQ�� �{�#���ͬ�	�j&eV+:.��]B� ��w�k �#�O��H�v�֧W�� �D����ɸ�Nch��"iC&� #�n�'m5i����Ɛ�Añ���b�D ;�B�}VJ�$��"��eb��1�&}�w8��S�[ i�,L��Vf�l��X�^`�M�o��P����o�_@��S��D��ߤy�Y���+\E?e�n����׫�l�.�
�>�b{�K��|<�K&k?]�c7%�[<�i�v��w)�~��+{��[��?�ܯ(�I����ɷf�`��Dj�4�[0�f� w3[�M-̫K�R��,ݥj	��gU5�t8R����Ci��*�������u�؏�o�����-��:v����e��Ư^"��'��x��!a���M]�ٌU�������Mb���<:�=/��Dt�KXT��~��E�L(��LK�D]�*�I ��V�T�����d��㼽�����գ�?Ac�L-�r��9n����e����h-�섎@0/)LïV5��[��&��rHe:�՟�U�F>U�,������k��XlxVHYEB    1041     4a0��f�K"�l�:3��-��g~����u ��8�F����?v���� ` $���t�agFg�WqI9��C�I��c��Y��t�ҫЙ�d�1�O��--rD	P''vц�M���4�a2"���qK�5�}�R>o�Ň�Z�w��/��ˉ]�7��;�{~sIE�7ל�^����2)��$l�=E���Ö��P��a?�x��Y��z^����K��! #ʀ�#�ʅ������#��m�!8Mĕ�GCD��CHtt��� jih��I<�dX��Fܟ���(��2 xH���L�C9��Uͤ
�r�c�ѳ��9�G�����;mmqIo0=]ե�@��Z��gdݍ�����_`O�|�Bu�4,�>�����v�ʠD�I���Ϧ#yTx٧*8�p �L#�M�}a���J%��<�W�[6VTP�8�,X��q$
��Z
��h���Tl��5��r��I������=�b�K[�U���.�������Ie�����$��������s�D6��]/J�"�iВ��2S� sF�u����V:��i�^�)ss�0_cC��_�k\7.���s���L9%0�.1w�íB@�����o}O�l�[,�G(���g�䥍S�8d�V^_:?ī[�)mB��'������d��Y�Zk`H)��kJ)�D�RZB�����*?�$��F�J
3���Y��ࣸ�MD	C��C��7��BT� $��^���Q���加�,��N�s=S������������?w�:�5]�S�|u��,@�Zk��jp/���(�!�:�2��{�Py��h����<��Kr4{�h�iW�j��ST�`ޮ��2��u�ذ�ț�=?��Z��i6t�^�����Ok/���w�j�9Vc$ព}(�l�&�
�!�V���
KIچ�UU=��\{I.�
��^dK+��a���������j�d�r�"��TE�x?��J���d�c�_�!��M53��s�B$�~n�H�l��˹v� �S��G�D�g��|X\~H�h�J��%O���p��I�=ˏ���j{��5iי�#i�2Sd:W_0"�������hY�E��8�X7���ƟAjy�Ź,���M5(p	Vg��ijq�����ه ͑}.GAѰ���{��ٟ(Wyq�XI��j