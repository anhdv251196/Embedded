XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��a���b��/�|����Ks\@�
��6� -@1�M�΃�����4��dM@���P��6�p��2�K��L'���	pC�9K�[�q��S�3]���{�h�� �G����vV�u���.yx��b`}����0't;��/��*Ƹ!u�%�d�r�дW�� �����=�%z-�:��e����c�[���6 �r������NF��%�E:+4=u�-��ȿ%��U��q"��g���k�,���{!&�N�¥�[�L��2h��f�hj��z��dQ��R�EB��(��Ȭ��u���RaQ�m�lp�3ctԁ1W�v'�	L�ȳ4�',/U "�T��x����Z5?�l�!�-��z�� o�5�Կ��"��ׂ:�-�F�iG �-C=�љo̵s��Lӯ{��A�ec� g�������]+�~$i���u������*=)�_P��nhx�(��E��_tv��Q �>�H�bF� �FF.�����:��a���`%p�����&�K_Gb�~-��5��|rɊJ��Y_ы2�9��Y%�{�~9a`�GU0Gw���y?�uzR�m'gR��l	�YP޿�l��BC�"���%���s�������I��.$؎�P%����Nl���Mc �Z���*���5�i�^�QR�C�Oz�GkE�չ��p*��$hk6�%a�-#�^����%fG@e���V_��b؁7t!��|���7R�� 8x� �9H	��m�L�D��FQ�5�����XlxVHYEB    1cf8     790(>ɝ��S�V�ӚZ;u%�D��}��~�?*3.O����V�~��,ݝ�kny�7�Y��@��f㘢:���Y�5���ͯG����b�G�N�x�w��I��,��g�@��`��� *^h�lA�CZy�I^�e�]���ŀ�4��Kᝏ��}�O,g��u���k�o���� v���ń����P�`�Z��awD�J2jl߇�b�2��]qli���_�V$<��_ކ��-��~�eJQ֊�>�Y��3Ŀ>r��S����#��;��M�0xl|���e]��'��y��?ބ��x�Y��	��$+����i�#�okBg�V�"�2��ŪbK�	l�!�Nu���aqH�pV�ը��=��՘i"e���}kI�o'f^���r��0ؼr|Y)���7�Hw���^�8S�.����ŭ�;qû1ǣК�k���fF}�ƛ[��ϲ�sS�6�Ԩ���ï���6��Ig��g�"�)qCtd�jV:�5kV�!������-Ƭ��G66��rQVR#i���$�(�Y�u���l�i"�4�i��]&mB�`w/z���h!UƠi!�G@�,�+��Ӯ�3��ݘ�J-hv��V�W�����sjC���{��;�ńmHi�:�p{�u�����w�-j�~�k#(K���a��Va^�Ɇ�7�Oƈ'�蟩|�]^J���%�i Ak���!�V��FxP��c�M��n����e�ǡe�ޘ}��n1s���/L�Q����Tb�,`���-G�<�Sx��7�+3�qZ|�Y������I�W�����a�7�"�/���y+�Akʇb�^-���B�0�]�;�H6���w�+X��͔�F�w���'J��'�Ig�g/�l>�j`bA�kf��4���
�$	����ѵ��TY�ݠ �!��B��1�Q�z/YY�>"��H�Q����Y��x��ƳV�&@�����������BQ:�	6:q�'��N��imC!��#���脌�<�":'�@�����s�p捩�Ǹ k���!DWS
�{`э�BcP��Cȋ"�Zx�s���W�'�	��ix%w>�%���A�Xv)���̊�������gi��=e�-%ù8�>�&QbՉZ�!e��lKy�s	2�J?b9Q�ќ2�v,��]6�Q�����H5K��=�d4Ӄg��Z;�-g�g���h{��!x�ݷ�dw��?h����vb�p)��H_l�M��4�%f�)8�����3��_o�앾ODڅ�����.��v,<U#R-�۪�?���M�;��ek�r$����D���Z�P�������I\M�`����|�4l?�� ���g���=���r��*��Vb��%���a��.E����_F�EŰzU���� 3B�Jc�M�k$Փ-�5e��x8H���p��| �x��{�O��E�iCk����u(a�����!�f���XNJ��Z�Я��υ�S��������֩q	U�5���Y�lAWYK�;���p�E�/�<.��) p��8�����w�d��M��$�J}������y:^��7}�2O?�ܟ�Α2�E.5��Eo>���#Ɲ7o'�W$qJ�6F�JD�CG )��Љ��!��M������
3�s��[�T�ہ��	мO�~�@��m��9{�%x���Z;�wPT�Gk&dh� ��4��<P���B=ܳ$�>V���a�W�S������cN�~��"y��ԽU/�!g�kY���K����%�i	u���p�o����/y� ���<5��2���pi�kfH_	o�Ň�Vy2�qOKd�i�ia���=��Sd�~^�C�-]��F�>��!⑶Xb�����ES�%�=|UF,�A�p��0�D��1	2���4�a�*�f+G�
��>W�-n�t�e���ɀ<�:��	�1y�5