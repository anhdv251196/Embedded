XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���
]�<�+̛bźǘ����Ig���I��p��~�f���C�����L�2Ho���y�<�jc��������:9�Ε��y?����:�)���������ܘ��ϥ+O��7��>�� H�n�*Է��-�r�ql���.õ�A-���Wm����Vg[��D����S���}l��~L%q�x5��{����_,����g"��)}����y��BtZ-����	U*�e���x�>�$��QT�p��^Wv�	���|hJ���8��Gh�C����G#��1�.��Fz��x]ږ�� W�ܢɣi\	\#dj��t�X6v��s� �0�Y��Jĸ�?I� 5w�S�*�2_�A{�[�J$��<�Z�Z��,���Nj!1��Y�)|���B�W�ze��ը��Y���;-ֽ��t ��4��e�Q	�?�% us����ঞt�`�^��u�:��륗�eu��.�.Um�m���lT�Ő��O�ׅd���n����c3>ݣ��@p/
�$|g%�X���S�}$���}*����mj����ϋ�֌����D2�~�e��[ZQ��х�h9�sr��'��-��4�ʸH�M��D��o�Dh�b��#eT}���tu���9�덖{<�%�B���DV>�Wp�p<-�t�r׸[�DG&Pr��
1'�K���t�-����iB��E�^��ղ�/�9 �]��J�yMn:e�J�U޷��)�7\���p`�C=ҏΖļ��Tv�D�@���C��N��XlxVHYEB    38f0     d30�З3p��r��O�I����O�.(��M�_%Z�^ՂH�!�x�
���S��ñ�\�#{Z��kQ4�I�[�ۃ�=�]WK{�u���D���"���ǎ�]�o���u.NY��(��3�>O��T]�|����PPҖE���6Gn���9�-�6�@�Jį�go���j>���8��7���3�偢A��$sh��H�-�nR'W���aFS�|�@��S�zy�,Ͷt�+���]*�!�Z�}���'g�r	�?�n�9��B��D3	l(��	jNi�_��?n����D�����_!-%��;)Xi1�YV����F�R����Wb��$M����?a������N�.+4&�ZS}u������du��/A���.A�N8��Y���V�Jx��B��%	���9�.�Jn-_��(L��l:��-:E)�,����@�	j �x�ڬ�H)9Ғ��Bi�7�5gp=���l4D��6Pj?�r��p�%���i��e�^��,L�T=��{�D��XE���v2p�SZ�;Y|����r*vg�0�
{Н�4Ї[߾�'�WW�e`G�@Q|���%�����Y��)���4��CN9:Q)�;P�vi�a���]�+�&����qs�qb�Ir�ȗO.u�c�	�@���6�ee� ��B��#(?�r���蘵��P��,��Y��W����b4�BϢّ���x�n�R�>���m+������,:�4{���	A�F��������1�x���IX{�نaY; ;Z:�I��('���Kش���۝��Ľ3�*�-Ջ$�<"�yi��"y��?B9�K��V���Y5k3�����L�|]7�	:R��!?"
C%��ME�YR*��T6��墐[�9xM���$Nz�0vMz�㫯ąF+BEP�n���}ޙf�fԋ���A֟˨�8�nq3H��p��v�8 x��Zk��8�M-߳l�CFӮu�
������v�D���rh>v)�.��dg���	L�U�4~����h�?W�J�ri	ӟm*���ڪ*��r��je�A����칽���"	o�ilލ��x��
9����x�}'3F�?-<
�����/oG;�Д[�y6R��� ��b��(l2P��u����|7瀢��|K华�c��_G;�ќ�Fei�m��K�V$��cr�_륙���ж�<�oiՉ
�<��"-*D�>�Blޓ<$?���H�
�C��;�C�a%O�������A!�����mTr{�~"Ԣ��	�~�4�>�(����X|�m�Jʪ���b��u�)RV�J�/���{Ba�z�N^�N·�N#}�FbI���]���z`=��`Dp�|����ザ[��Z��$�kw��OB>T{��y�κx>�íP	:~���i]8�� W���I����0�/����Ԓa��G�i��\7�v�p�VТ_Y�ֳ�����V~�rI�G��4�y�u29�͛6�D����5*�����l��2�
�Ur�����h2�v�M�`x��=��q�PQ�@�e*eÕ�[R�2�a��Nw�$<G���`(�����P�+ z6�hC�k*�U��J��$����� ��^L�����'�砂'�����nǬ:�zT0*9��T���W6��-��+��3�@U���ƍ��n��C�QKe���xAM7%E�S�E�4/�e4�=��A���t�l��]�`]�ed{�N�B���0�T"a�|���PNO���p+���U{]�Gc�Զ�䀝~����	R���[+(�yWKׯ�e!����>O)�Q)7i��m� �-H�`�������ie�/W�s;b�	{'�7��B�֪�GA�f�N�����7o�#x���3t#nV�5���	f��)�ETz�?[��+2�;)e��W�v:n�;���K{<�iKL*���"�'�y���ϝ�Y8���0�:�b~�����L ��ȉ�V�6 �h��l��s�k���8���I�����Gȸ��m}���O9�M�{� ��"�|�na�.��/����ˡp���|MvG��G����ГƦe�@p��=�M�W�Z�#8$�n�̷,�&]��n5M���O=_�J�(03<}�}������0ȓ�BU�&�M�;���� �d���1n9�׫CQ�QR�A�I���	+��N���k�����D���]����h�t���k��|
0x�eJ�0� @A�,���N8��)�Ǆ8pEb%��0��w�Ky_:�-d��O���ى�C�����.�M��GA:`;������{��Qm��o/�,��M��=`�?r�9&��\�G���m���]s_����kU6���k���7��2�l �"h��s���E�����&�����"I4�ZY�ea��W'>���(�Y�@�p��рulp0KKn��¯%i|�m2h������2�W����r���$��ݿ >��]O�K��ep%�:0����w�E���]�w`�T���㤁�!5.���|���$]&j+Qq��Z-���]v����<&j�Vl�	�Ŷ��=8��I1��}��pΰp�:-��bnr�c�P�7W-��*a�g!k����y��g��avhD�"��^�= ��d4�d���w3+�^Ľ���G���G���g�AY~�̑��S�׫�2��nʊ��R�-����R{��ʢ+�m�5x+��N���J����;��^�.��iU�l��z�;h&����^nq`8���C���U�+��-0���<�-�������j�^
��r�J2���vE]��&R�6��cWWd���k@���8�c�J���2$�:g�?F&���M4B��ͽf�}#U�i��۔�z�9�}Wj>hpb.u/��)�p����p+��I��'�$�ߦ;Km|&���-MR	e~>8x��߼ ҉<����0W��PM�/��*{�sၙ7���{
���Q5�B1n�ٸ����^��K����.�B+���@S���x����ic��	���g�t/1j��Jũx�F��$џ$f�K�i�_������80�'O�;�jM{I�\_)'���b^�]&���*�bi�<Z�s���y5ϒA!h,�ų�c%���N*c����.;�i�}�Rg'�g�j�x/��}��b_g�5�8�<��V��|���=�۾Id�Asd2t{W�yK�\2Kd��"������Dd"�S�0�|��Z���Ok���R���3���܉2�f�,?��f�"��(S��v��7Tt�5�v��w�m#�����pc�����