XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Ӽ��0�s��o/p���]�%�g�
+��sƸ6'��z�^s3^W#U�ge�+��Ucn��>ϊܴ���;�E����؁Rc���>����P5t���.{d��k<B�0�����pW��E�B��~i��粑h8�����dg�jD��u6a��R�.���y���U�-���ď���N��Ĩ5��ՠ�X�H�"zGI�%���R9�m�ʈol��_@�$��W1��~�'��G�������Av6�N /�Paܲ	�Ϝ(�N_t�����p��맘k�b���7R�С4z�.�ٽ�����Z�>���7���������腦�(f�a��Y�ϧ��Mz��2��#K�J��u�X�p�BZ.�H���o��(d��%;h�m
�d�Ғrg�ۄ�&���أ8p�������.W����Q{ύ��'Z����q��	e�zU���,!����$;?���$:p0���w���!�|6G�ٗrM6����I;Ɓ�l�.����p(6�oULU4're���vsT���R���D)L\�$�.��۷}�lڞ�7�ۉrm� ��zy�m�ow��V����L	.A�P^X�Cs�O�������?Xp��Kh�3ܖ�ɪ9���[3��9
�eH��
�C&Y���;�Qq 4�9��-��"�xգ��4;u�����	@a� ����h�4�8��OV,�f�M<��/�1�*�T�i��E����FY�ɄSܪq�����H3�v�;��ӆka�| �XlxVHYEB    5ff4    1040-&a�?�����{V�N��F��ae���u�02 #(���)�S�$��<nE��إ����ˌ`8t��'�i���:o�.�'!%�=_�˔��h�����͉]T�+����IX�b�es�Z�������!ǰ!��E�9���F�^Bj���u)�����X��MlH�|�$w�В�ѷ�&Hye��ᛀ���5@�1R���PsL�����1B��I�F��[¯�JK�uC��
H_mlä�`��"	Q��e����+�S���-v.�":X�����y���ڭ�Ĺ٧*?���%�C����4"��Ww����/��J`�c���o�^Uj���x��n�V�a�z-vu�-Ks��>��Q�T7�R4���qSo��O�c���t#12ll�a;I���.�����c(��,W��o���{�C'��ng��qc�������*��N��;ix"��WB7�A��~2#Wm����Rʓ��3�ﭰ��m0����9��CGtG��zL��J�C��Z��1�[��C���Lp{�4�5��Fc�xZw��ĸ�K*N����a'C�~�\8Sr�K��"t�ÝK�l]�e������Q�o�Ɛ�t�Qea2�?_�K�$GV�۾���1�a�8G��	H��Fв����h�	�c�ǚs^��"�_�B�z����C�������{�Mq���&�8p��̝oD����N�S� �Bv��`9�y�ޛ�	��`�ZHO��v#�*}�S��S�"�+C��������|_���BK��om1��5ɬ�`�x�Є�5�g����_��a���;�@f�>��:��s������#��vi��7H%���Υ3���'�%�~-�SEF/DQ�o]�F�~i֩�2��|����������2�/XB�B%q`\H���lϘ8�U��K+��+C'�ܣ�b�BTp��cV ܿ*|��Ś� "�^w�HlKe�)�uj.)���h;I�Gf��&}��f���L�O���!:���È�~-)����z�=nPmp�CDۂ.bd4�ѻ��4 �7#4�A.7h������K�5?�{o�k\�!��}�S#v�@D=�؉8&p�N�Ni����D���K�E�ۧ �-D��Y�>�e���N�/gύ"�0�iG.(�`�ۊd�p�>�mN�pPH��:0|:��N����F���қ���AD}?��d�=c�.̪ZeU��Ɠ��ɜ�0�cRJM\���x>��z��K��^�y$iT7T��}�v ��gh	y���^N'��U�cs�9|����qz	��Ihˏ;#�%�<������=�)���IS1�Ǝ��@yr�´�qbrV�ZC�����kyG�(��1�&ǥOSG�U�y�k	�7y�e�I���l�WJ(*,Q9��?�^�zH�l�!�h�x���&�C��/_��<bG�e��0�9��F�y�o�dQPF�����E��tC��S�P&��G�yq������wHN����öW-j����HrN�<v�鄻�U���h!��S��N�p�B?��{9>2(_��3r���3��ͱ�E~{�,����۴;8*>��Bq�c����z;[ճl)FUoT�H�Bq�L������mPf@ϪE��&��6��!�+p� ��d�yeo�_���'	h���$S�ȎZǡ�~O'���C��9����� �_TӦɒX��?�=V����`=���9�K�$o����~m��[q6fI7��Q8n�?���?�(+ņ��϶'���0}��J���
^1_˸i8�d�0�%�p�
[<A���}���;P���k�;04�?/p�@=3��Z#�9*�8F~C�r�����ι���ؑM�N[ɰ��6�Wv��U����%i��uۖ)ۣ��_2ܐ��=�����:�G����MpqF��0N��`04YC�"��4j���jj`���HG9C�/�y�dy?Ӿ�Ya��(�=�]��K���&EsrKtw�Ĕh�SF�%)���;K:[m C��]i�[?�ݙ�>�+���9���x�ŀ������U��-C�ݡ��}�Z��^+�{���	���~�˭4H���C��[&���� �e\���S�ΞPg~���.�ʀ�ih��i�F�A(%D��\��0����� ��ias Vv�P�i��~�Gﻟ�>�n�d|��$��rT��^�S�D3s�"��Z׼�G�9�M��֩��S�U�I�\�?��9�X��Ɇ�%���e!��ܘ�����YD/a���G	Gψ��n��<����e��1�����J�X��0`��'��0��	
Z�F�>N���G��\ٟ����-l�H�ڜ��?� ���`�7<�S�wd�b)i>��Ϲ�~���Ms�Q��d�U5(�����KG�i��d�s�ˆ��h���s��@!�Qׂ�k�����@eqkk�0�"f�9�$���	��*�c�_jx����P`�ے�R�م&x�O
�	ηK�r� N�qP<[]$n"~K�H�vB������x�f�t̷D'�on�+qp $A���܊y���g7��z�֛�[�k5����,��W�(���~������a�Z<�8&Yc��GM"o-��p�7����m|RBŜ-j���Y�ӯ�[@e5�ק۶\\M>ǓRQ�h�0������c���X��CF� f�|����ފ�^y��t:7c���o���2 �b�֕�a���|еb�%�>�A�I��.i������f�W'ʦ���^�JMa7_�ǯЛ-�s����o��3�����3�c�M�.���
��X�
��ш�y�����M�+/�	%�7����C/vH�'��0K�1��+^Z
c��k+�Eж��g�_H��+BY���"u���ܾi�v�^ݫ�[K	�U��S�Bi\`��v�����b�~����������
3���T꧊MW�#,�m��yP�&�Q�GA=�[�}�"�:��u��`jֆ�2�ށ�982�f�+�9��VJ�Ǽ|NH�����9d[����Èz�+t�1.�\*�����TC�N�/q�dd��������"���2O@�¡��mCߜZ��c���oHzTI�`��5��
Oo��&�Uv�J?�Y����r�G���h����1�#%�����۔u�k��N��!1��퇋�*��_T�j�y����^Y_����+նe�9�pКVhS�|iM���&�n��<��Sh&~F��U&��܏�u�e�]�q Z�u.[2%�9c<�J���͖OUH�|�s�2��1v%����>q�w{�b穼SXS��톨v��t����^k�z[@�x�P�ٝ��1'{Gp��O��E� �U�_�Ϻ��`��2#��t�H��)Id���f�$Un]�
w,�N��u�j���]��ܸ۳��/䰖n8h�:��HI,�z�Z����YF�>8�޷�u��?��R�$�*p��|���]b��iJ�H��^��0�]q�:r�ϳ��e]"8���s|c��ţbVR	�w0�����N9���ep�q���XL6Yr/{c/��9��67Z���3U{���	l<s9�)tL�#�n�5�>�'��K�b雎�=�\a.�ܯ-��*{w>�Կ�o��u������]u����ڛ��;U�	 ȩ�M�ר�/��v����s�]M�%MM��5�cKtW��3!��uGnc�<��5) ��4��1�K��/�`Y���y��c8������U�;�G+r=����;�����&~�7I���ď�+A�ԥ�s�ʽXG��w�n�`��x���tF�����6ݗ��R�omiDz��c��/����Vvj��m��=��@ D/��Nn��8�� R�k��g�${aO�) � ��%�U;�Rx�p$!jW.��	�7en�`~��Hr��V�]!���ڳ��fz�ۭ�l~�ea�Ѫ4�aG�4@B�E�roĬ?2q�X�G�\������K�;���\mx��I�]��f��������l�Pz�-�t�0�͛�x��й5�g8݋ni�YgS�1ڮR�b��s�a\1\1�Rl��Fu��Ό�_��%�I,��