XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���Q�D��X�L�eL�FZ�Z1�2�)#�� ��F���:ݘ��$($~�_uwWI��l�ī�퀢-�~W�Tk�<q��;��?�(��&��g�z*e�Y���� �t����G���"{*z#>C9�/�h��׸�4ݳ��;-+�u
����싐/v`RA��6�ld�'i�[~�fW0	
��XUO<'�!j�{1&m���ܝ�?���S�f�L����b1�yU�'�[o��n��F! N���H�&�꽻爞����xi��>��i���]U�!Po��o��� �Y{��mP%�mgAo*]�-��RF����C(䲩���:b����j�v��V|��R���y���]���ij�w�Wk�ÚuLy������C��nY�^A�v�|��z1�-�ܚbv%�-/��A����?�$}���s���:'�qG��UB*%�T*�y�ӿS����; In��E���U�hauޟ��Cf�h�U���#BE�=N�z.l�ĈΥn0�M���g ���#m�Y>�N�Ig��%vL�쏑QO�.:,�2����&ɍ��-M:IV���-(�؃�IR�_e&⭢�Q�H~���fO�J�>�����(�3WᡶFyz��a VU��'@�Q��\G�����Շ�E�����u/d�x����M\���n堸�Ŵ	��F��ֳ��a��W�k�����侧� pLԙ��j�.:�}�Yl=�~߇v}����嫮d@� }W����,5�]�XlxVHYEB    fa00    19d0���.|����P�'ظ<�o�!U�S=Ӡ���CGI�J����k.���@��E[����1�c6�=�#�	��(�ˌ���nA��Kq.���Ƨ��GG�p#�եT�)�b*`�T�Y�I�خq
��v:yl�Ea��j�9�U��;��R@2R���Ş���]<A����}�dm �7A�9@#����ܑ�w"P��\��A~��.�wgd���U�%������-n�uBbkv�Y��E~��`���+@��;�`/+�U��yl8j�%w�2���L�͋c�J��V��3�z
X٦�w�g�w�K�>���Ɠ�Uz�P��,J<~��w�\�t�X��k��;q�͐v+|]��ӏ�P���{r\i���/�s�\;=1@�,#ge�C��vM4�ɼ*�N��Q~�:,|�N�ۡF�E]5"�l�y��=�K�ȩ?	b� )���[��Ҝwsb
�QR���~=�L���\K=Js?�N��S	��ָ��aF�nZ�D���`�xY�r�ٱh!��(R-řZ�=Cu�u��=@�;�iY2�]�ҫ�nd9�� :2��vcM��7z~We�.���͵�����4x� f��H�l}*鏭�(�'��!�1.5@M;��*A�J :�]��9m���]o�K��������
lӦaΊh���3)�U<M`Ԙ�`�����j���qP�uy�d�f�j,�o�\h�8�?�c�G�c�t��k��j��SA�I �jx��������Q��{2z?ď��h�����.��%��pF[�����u�o���2(�q�ڲ��W����� �8Hb��-ܰ�F��7�����b�M�d6?�d���1�*�'U��C�B�x�x!�I#Oi�+{�y��V�X`�Q'� +�s���Ů�G�ϯs���d�Lt*>4:W��Ji-�C7��S;��1�eC|�x�m�w���?Yq��prw���G+��KQF}#��i�Ҭrv�ui}�9��y`L mQ�+dM�
'1���)�y�
m�h�g���a*��q�	�(�rK�H������%W�QI����"؁n�ar0QIѿ�0�s���������6%�|�y��)��cLY�� ��������@˿I�<o�:�y�]ٝy�X]��Ř�Z|�4ہd��;U|��+\ؘ���PT;��d�퍀��F7Y�3�^ ʠ�]} {a.�M#�o5�p��r�vh����\�6vwO��-��ڻʐ�3WX�ur`�ŧ���c�����Rq��o��nQ���_�/�du �X��oT�x�^���z=	�{� E�� ,W��O,$8���!�R��I�15�RŠ���ֵ��G��ߍB�$�N3����k�K-V��}�#���Y�OuU�z��T���O�u�Br*�tt"G��O���Ԉ�R%jL��:q�e_ݨ?b��?Ku3��C��?k��"F�ƭ$1��.3!�"�P!Ւm�yw��$}��HZ��" ��_����|S�Qa�\��i@��N�R:ב6c!�#�f*C.im��>�_��l�,n0ՍVf*��]H��i6�`T��)�S���*-�����F ��ٹ�Qt,��p����gӝ��z!��u2�Q���dk��m�2�/=t k&В<������G1O����"��OzY��<�ѽ��LiM�=��jnI��� s>DbW��ȁ�{��y�9-���C�o;|3ƉEy����2me��>��¨��j�%s�?E���%~����@�)��K��A�
�L�ؔ,w��X�5Q�:@��<�m�N�z�e�)�+Pfn�lw��;�.@]��pSW����R_�3{�/i�(��n�࣯���Q ��3,
`����?�E���nu=j�	�f�4�^$��l��$ ����%@�8@�-(���tD�H����iro%?�Գ�%�fTH��@4�T����y�~��qӗҕU��"g/ l��;@=����h�P���	 M��%�2O�8����� Ͷ�͇���t��H��!�\jt��T,!,�p��Ul�#�X?b��.�I�~�c��h�ߊA�SoK��<?n��+A��ҡ�>.�*3Y���6p������B1�CR�6��g���f�DɁ8��25���Ft1���g�!Co�T�m��l�|2�e��k�$�1 ts�8L7���+A�Z`i4��}�r8�+ ����	r��2!�|�F"Gڸyΰ	浪�f�tVJ&r9v���t����� ��3�F��*Tud×kC�l1�o�U�K{�qY��ff�ĝ�;��{���Y�yo��Q�_��4�@-���� E�)�9����*����ݾ�mS�_ =]����#��&U,�5�8(�[`�,�S��'�k187f�d�x�H�qƵ��'���Mg
��>�V+vg!�����R͠+��������6D��;�4�02�^@eTF�[��36
�7�B��K8C�ّ�)|y�q�-�m�A��;M��r�)� o�R&���B�]�,�P&S;�[fc!X�$�S��(Ƴ��_�I>���!�`p�K�	E����1D�+�u�T~��B�{����3|����|8���U��%a[��0��~r�+�Mg�f3�o'�ƙv�A��f�9(Z%l�����Y���ܘYQ�k�R��<kȷC�#{�h�0�=ΐ4����]����M���vnX�xSh�`i�"��M��/Lg�7b�������Tq��Օ�1 �Q�X��F��
�C6|Γx2
řB���ýRA�	pl�n���9�����$~*��r($�r��AM?�Ҵu��.�B�WhbY7���&VĚ��5���<��91�b���m��K���:'C��P��gj���l_��mPn�|������w7vAQ�X�f���{9��}�� �<�2�>\�W�/�z�߆���.1h5���5�3��T��.�_�P�LVtNfrZ�0�aHw�<F��v�"4H�P��J[�({��k�5?��gYda�*7�4����Z��=DR�ۢa���|�ݐ�+t���VZ�7�Y<�q�f��͜�܍]"gI³7F& \+��:sjOo�o�fYO�%�!}��܀�p�!�����഼-e��ð�amHg���v��,f��{�к���ͽ#��mPt��m���(��;�U�Ɨ�?����+����,���(�t34��� �����Ck�-n$P��	첬��M��}Iz	�()\=�U5?�����LO�7��܆_Rw؂���Cѩ��ª�c��ў���<��"�1�Pﴲ�gf�2��!���A8����V��w���t��! Y�w��͡T>x1�p�\R��s��H����|����u�&�eF�sv�͂�v/-.�zO�4�v�v�q���~ dw�@;2�*��]^iZ=8A8�U�z?b@ޛ��(/F4��X������ɒ��Ї���Ab�.
��,(�t[�C�h�-�E���W�ׁ�pz�6����<�A�K:�O���c�a�A���͍,��OYFFZ�o^n��Ҭ��ڑr�7FPI��'��f�2t�5 ��Zx�WQlU%�%b�w��S���L�j�S��/�g1��f�p�%��d��J�&�o�H|�X#%���[$��,"��][�ʾ�v@�0�q5�'��~z��PAx� _�]R	A<�������k��¦�]^����H��R'�~�"@墟�:�X=}Ne�v���-M������W����N>YHGX bɴ9�:?��M����1�6	���})-�}�$(`�P^��9��T�dwRE2��3"���r!���XǶ�cϤ���F�NH?�:2�B��M�(Qծ9 �5�S�H��u  � ��ڌ3��/~O�=��D�[�M�I Q�apQ�Zb��<��t���L7�8�+̾؋b9��8���!�-�vo�a[;��=��=��R�3?J�B�\vad�A�@;m�1~�O[���>U����<��mw�)c��s�\�Y�C�M̱���1��U8%�ɫ-��m�]��Q~{~/��!b�GCP`���]�A_ɖi���2��L�p�Jq�S/A�W�6�9�h1�!�#�2P�TE�d*�q�.g�d��A�iL���Lf�|ÍAri���z�_�ٟS�K�U������0�>���|<�J.4Q
���eӅ�;b{�I�y�[U�T���px���3I+�c��1�unA�\;b�>+S��Hm*c������yd���v$���1K_�s$�2�O�: �/��o<�{�D�򑹷�Se� �V����/c���)�)蒐�ҵ��e�0] 㕎Y��a"p�����ԦCc���'2��(���3X��l[~jq�#��8�������"��� ������^��)�z=���%��i�a��Ds6�hϑuʸb�i*[G@�����z���U��ĩ����wm�(y�����he�\s��mڅg�ҕ�6�u������toʧ3?�2�+B��22�h!̓.���,����J��fU�.		0����rA����:��A^�xre�c ���z �i����˖���q��p[U�ASm�t�6S����L<SRH�y�I4E�ic=�k$����W.K��f��1�,;rn�E��\
�e4��;���)1Q2�0��v�9��N@���p(j�n@g���e���9"������޽��3����{��)Io͵�	��w�0,C?�����5?��o*VC�I�'33G���E6�Y�[^�~��6=�o8)y�\3-q��R�qR���uN�3H�G�KƱ�S�\6��.��t����~^�������^x��Z
��ݚJ��v��ڽPŵ�G��isCW�4�ң�'Y�����,!���k�#�Ä�3��;S\sd5�k��NJ�'�-��\.�:�;
hUh�a�Н��$���(�3B������y�u>�H����¦&o���8�0a�j���:�������UR�sNP��v8��7�C�l���8)��J��,ޫ|�J�<ϳ"a�D�c��L���Y�g��2 �'�S>��y���K+0�/ȗ�Y|IlO2�Oӿ)c��!�L,9
l�tyqעC��xG��	(���ץ��ϦQRT�?G�E�	,R!��ÞQ���bV��{[�\R�Ӊ;6�nE|Oʮ�h-p�Ai`zåT����]n��n���4<I*u1bE���V%~����c�� �A���V�A�����=�e�O��_A����M��nF�X�ض�04'㰈|��z���Y_��^`�u��Lc/�@�$����$�if�-��p,�$Ev�����]��#c���T�H�.�dpmsw��B���q���.���܌�£��$e:�L�RYr� &��!N�R�L����VظٰbГ���9f�0g�m[�c����M��g��6P�w:@w߭���l5��B��m�m���W�^;(�!$�ǝ��>VD�؂�sU�a���;�ˡd��	�y<�a�i��=J�W�Bͣ/��������#k/<����Sd�/�cH�41��)�K���ژG���Vs�_������]���|ۿp�!�G4Ɖ�?�ŭ�8m��,5� �|�8�|T|��J!Z1�/��z{2~_�B��9"�1SF���OT��X��}���ȕ8
k	�J)b�#����+DZ�>��|��W�rA�-�c�`��N��.22���� ��]���/�d8���8�v#�{�pߙt�N�g�{���[�</�8��E���d6�1��)��׵h	~��v"Y�M�-E,�wFܕ�H��i��,D�~�>H��ժg�s�� 1+���F�0�o�^��SD��h0Ջm������4[K�b�{\���j�I��IVٗQv��ge���|�����mrN-n��FI��s� ���.��}�5qAk�1M�w�7+��6�x(
v�uԣ���Ϸ+|i6�Z�˃��}=�3�D�T��6��겔��v�~VFf�W�?(�S}�������  ���㏎T^/����P��̥Їb��'�� ����ŧ�Vڂ�4U���U�mn�[�ֈ�С^sM	�L{�gdMyW{A���:��!�H&�<�tg§�rJ�3��i���f���ѭ^�)�-�fX�\+����|����]����L��$V�ʊ��h��Q%���Bv�>鐝�t�k!O7� 
hD����2������+���]F
x��죔�{dy���4Y�=�\q�$�����6О�w�K���]�b�=�8�8(d��� �����M%��b��ǚ��d����&b.
�������F5�0[�Q�5̼�9���=���S�H�R*n8����'�������C)M����0a]��(�8-��x:Ƅ�[�Yz�)�C�b�^C�x^��g��5#�N8Y��9�uvAy��i+#?��xE}2�i�*IIt�}�J���>�� �.�{u�Lvc`NH�]))�Q�R��t@�2�xQs/ߜ�9�c�ή\�XlxVHYEB    fa00    1630��B�~�|����x�h�nJ���]o�k��>��B���&��ȥ��1��/!�z`�P��?���.�7:���?�bN9�y��`�6n�~��g9{^�?�U;��I{����<���%#��\e�s�.�E���w�{�RQgHS~h�
�-MXcH�����ԝ�[-������x���� ���_� 7��_#Z�!�R��a���NV�܌!���CzE�v�`\w��m�ܸv��[�]͊�:>|J�m�B±��
ͧ��d!����4�8'̠5LMĞt[�^d��TGA�����A��'�Ì�by1&�a0�A�j�N��#��Di
ɵ�a}��8%�)̢_�������b�$@<-�������8R�����R�VÖ��|S0�O	�S��k���CH�M�����x��0�&�����^�$TA'�qA`g?6�4m|&5N�;kͪ��Th�#��C;���w3ކ���'|Nkj�IGP��j<����/��ݸ)���c�����[!ʛ+�\��;lC�1%$��/!u� |׭�W�.����D��u�F��P� w*���K\��PS�[Q�˩~��}˝��a���y��U�	1��d:3
�yy�Z� o�k"z�	emҘ5��-�-p�3�oH
������Y�6ٖV��4���}�1�Z��4Wf��o��/4Q"-����dBB��,�Տ��f�Y ��t*�ѱ�Ap=��9qh3^�rs�`���*О��V�9!��߆�,��H�����W������'F4���[�d���a�ch9�� �r���AVp"�
��g�5֔��>S�3j��Kt7��=���V��JԵ����#�S#|�� }F���R3��v�*�+��=%-�Z��(�D�x����_@x�`�:��W�1���LE�T�m�X;H}��199��o��_J�Fo�x�y&�(��� ���X��Zh�l0e2ȁ���8s�pQ��Z��Q
�_)7#%�����"�]�d��c20!Ų�ٛ?���ٱ��/�5���la��o���ӎg;Cf/��02�=�kך��8X�e3�>��|DP9����5
 Z�Z@�7V�Jԅ�k���*^y(�:�4�h���=�Y�vY�ڀT ����Y�})?GG�A�[�S*�"��X/i�#�){��c�����_pO`2Q�U@�Y:��e�)��a)��)��0ׂ��k�9��KP��;�))g�OU��$���|�՛Xi�'��?A#�?'"/Oq�ž��
�LW8�"�-¿tz�=�ݰұ^�\��\M�Qڕ��B�!$rf϶�E��@R�����^�=$��C���P�I)�g_icvC㱫���T|�$"��+�=��n��.S��\yZ�u^/W\�ڗpt_�B2���0�� 6Ta~
�>�)�4گ8/���M��#.H���TL��A�iI�238j"!�(j�W��H��A!�HÑF��&M��Z]��2ȶ#%=|��L�<1�f$��#?zSm+�+Y�]yv*��7U����Nv�'�5x�Z��{�cQ{�S�3�f�t��h"/���h�;�F��ô+)~Ż�J�Q�:��zJ5�I7g?�gL&�P����抝�p��ee���Ȏ�e���x�I��m0�yo�?5+`�Ǧ`::vf�p<�vo(����w$-��q���o)�(���T��A�e��$�p��ƅ�����?�F� ���{���j�f�H�w��B�8�'�!
�,N	:�a3,M�b����ߩsN�6ah����ƅiNw�����ѫ��H�f��t��.��d?��H�n�����)�uL��)���\&f�����>dr�`Ɛ��oG���t�=7/ϔY�0��NN9�v���k������a���Os��Ӓ����X(}H�����3*�x��5h@a��Y��8[@F(d�X3�O��E�G*��5��\9�v�F�o����1nǸA����[�ϒ�y���;�YpM�@� �L< 8&�w:��TS�+��#�y���n_��h��	��6c��a�o �%���QU��7��^��!,��2��`�UOo�	��F�� ��x�N�~�@Ewα;�S��x�v�a�E���_0Fʛ�Hx���e)��˛�����(M&g�1e�H-x;�Og��~��8��s@�XB*p6���7�������`8���A�ngPI<�F ������Z[�j!8���Jn)���Jm1}Z%{���8W��M�{	�T>&�YF�lA�δ��=��B1�o����9='2�R����zAq�����K��VX�A7ӂ>ZivJc��fb�oz#���6���������q�%�猈<
��W7�i����p�m���ׄ �q;c�n,iDR��q�Cj�~��Bl/��:r�y@u�O�'�ڂ�vl��&/�#�� ʂ�&�q8��d�Ad�pZ%�;�EϹ�;ƫІ��l��,������L!�����)�k��3�2�B��W˽��g^j�B��=5�sl�	��Ϫ��D&9�:O�~���xc��ڈ�Ǡ���䑁7�)3>� T=��Ҵkvm�3I�,��\
*f�e������B�혢��ʨ�� U��t^3��:�T�����r2/�P���
�^�n�Fۮ��>����^�T����!��+�oi�G�	�w�@�EU���ߒeZN �&/.]���ExVV��9M��ƿ��7��h���Q`�e���?������񱄴U�ڌ����#��4j�WC�2�y�^q���HZ����ٶE;cw?�'��S��1�,w�{G;y��Po�<o����P�+H�
Y�1�^��˧@Uwd<�"�ֱ���[B��E�/���� ��>*X/��A}�?1�������5lXG�JY����5���_|�$"�:&��s[�rA쓣�r��)��Zy�/�mW�+��Bؤo��4�<��9��� P���i+��q	1�)�i�I�?�-�Fw,��6���c�R�oL4ˈ�( �,q�x�/ AE��;�9(K\ڊ���5�qߌ�.���R]�iX�o�Cy�u�'���P�0y~��B'��*��� ���>�t�A�G]�c]���S{B�Z�k$Z٭�\�HdT�Iր~�v�GDǇZ�9<���T�m��UQL�''	�.i��H�.�4�!c>8��r�3|@�}2�aq�\�<�B����[���UCT�!��`����մ{o�ӺKy�Y�R�$���T��bZ��N�s����RlM/qg��zAN��+|���7��p^���A���%B3����M�����V%��+R�5֕%���
��B|n~��_��0dJH�f݃8�{���,��O�)���?nu缻#�
��>�7�?Zg��A�6�������:�o ��N�[zI����P�9�o�g(ݯ`�6��?��8����~���xM�T-��}�NĔ��=_V��D�n:LR�Zہ| [�8%�$p;zQ�}�ރh��b���XpU��f�$�B�R�'�l2�p�LM��my¿�G���[���#��,�[��"�y$B���(��K���-����|>���N�r���!Je���6�_��~T-��C��2C���x��[�E-v�Q~�j��6bE�2Q��lW�g"_;��*�/ػ�y8����S��ik�$���B��Nk��'���d�#)�`�ZB����5��|�����_���5�C-z:�>�_{L.w�59~���"W�Ɖib�<����)Bſ���lc�l-��5+���]`j";K��|f�2{u� f^�S[���� �m��%\�!\B}%/�s⍿�\s}X�\���!\�����ӗ+��j����kǮ�!�{��g���M��8(��e2�T�����5d�s6N�_�O�ѯ,�2Z.sf*���D�/3�@/��`���:M��,v�P���w������c����d�Ű�E	�Ӄ f�,�Le��갠�/�o��yr���yj��Kw�ς���NJ_�T��HB��,��,��������p<r�K(�̎���H�V`�\��v�=g�l�I�4���#��Qp�����YG<����g[����o�9���͕ߌx���AOg��aR��c��L�����r[�U�@��i�	�׀�M9�c�����yۓCxV���L�OThS���_z�Z{U��ܭ=���+��0Ϛ�25�ƒL�s$��^�"�ǋ���;|�0>ӕ���>W*F�����>�~6��<��y%�-�]����g�{D�	X/���*�C�À(� ��b��oGg>z�?���N@n7�m�;�����7��"�p�,�+�)�)c]������f�]��
��!|f8��͐���|���ez�;+�y�1��#�*j��Fw�	[��t�AhX��
��1{�V���F��ZM;O�(Bž���hv�E5B`��%]�Q�v�:�j�M$~��w�M9v��@D/���:Ni�!9G!��;��n����'7��?�4<_�o��X�
+H>_RW6e��3�2�$1���ǎ{d_~r��V7����fz�A�W�x�������G����C�C�w�3�K
��(��6�qZ�������覮J���۶ˮ��S��z�/��w�XJ~�#U!�Q��XA�d��up��n����	����s�	������ϭc�V�/(Y��[�����)
�>ofq�N*��$"�=�t|��Z��<��U�
�&�g�cP5ñ�/�x�u�&�Ba8�$[]�a�+\K�aoap+$����ZD�ӹ.�ϝN:آ������2�4+M~^��!�����c^�..G�pT{���ՠ'3@%J����j��;z/!LP��d7�h�8cb5i>e Ϫ5�+~��un�+�(o�
$����`_b�g�u��.�Ҩ��>"V�(��Ca�'�h��*��}�V����MϐD�����wV���������0.��W<A�x�p�?��_�,1�%l�=�А߮@�(#:ۜ3�Xn���B���o��dt�l2���]}T����9�ϼџ��oǾ�]|�l���Q��-o��ߨφtr����)O����$���B�m����ۀO�F�g���^M�N�gM����W%���Ζs*��= T���a���ׂ����*��(;zَ��u3��QI����m���Nj"�:�����{̥� 5H�7 �k��Q	������<����ٻg��Z�οs�����u#�Թ�WrO'{^�uuѷQ�yǔ�����&������2��>g��2�bN��@;��}�-���-y4mcf�-x��V\x������F�K�I����4�wT��
�΅�"���D0���^�&�v=�֑�KJ��*ߩ���F\�����ٛ�I&,c�{��I��ǟ�!��X/�A�A!����o��㖖2�?Ă4:=��u�}�ݮ�XFt��p%�����`���������}p�?�1�zk�Q�;�H��m�\��Ӽ�]�7��'ȬA�e�Q�}�O�;Fd���­2h_G��͒�d���H<��/���#�3����2�X�O��:�qAL[��XlxVHYEB    fa00    16a0��k�	�?	i�ԘrVn�K"�P��bKX79�<�*�D�;���J�)whh4���K(�?~���W#�<"2�<+�%�f\q�K��[݇�|t�s��@?���ӽ=�}�Fp5xZ�|4!�\���p.r�?qI���5v�C8o	����	D�������f»:�2�)��˖)��&�@�ե�q\rM&k��~���\�mFF���9�d&����l���)2���/r���}�*�ZD��n�+��m!!�7X���.�aF���,���4#�uL6��L�@euY1�Q)�pαi��"}E�A��wfD�C`*�5��^�#�#/���"��q�fP!!�����t��d'�TF(�D95d�k;$*[��W���맴��<܁p��vx��3}��KeXm8��>xbi�[��~+�6��G�*�!+�K�ف�Ҝj�o8���j;��sȤ2U*>޺:��M�1"�n�(���&��z��.���ݺ��Tȥ՞�X
��� �EeK'3h5V���׫�^�m�U1��x�]�%�}v�)q!��>T<Lg8����N�E="�5���2F(r��kI���M3����>�Nya^K�_ʻ��Q�m%��yf(�17�^C�s�vu��+��y*|�c���1��"+JFF�?�`�΃�M��S2�E�����z�"�w�L<mD��@1%8�����r5�5�O����#b밥
�\D5E��Mjf�gT�Sd�82������1Xu��21Nq흷FIq����w�[���M`��� �5��,�v��F�}7��ʫ��>��<����}@��8�A �F_H�7�H#����lYR�P�l�L1�l~X㞋�{��_Ԑ-ȴ�c��P��=�.�#��ݗB���bR�JR�%�����ǃ��R`�tz~ҹ������������q����>u�o����ek��nbN�y2Hɰ������k����e����|Vp�3 匈�o[� �I���Y�\�j��uKٽ��-��|���[ )�ijAf%*� Ԛk��lQ� ���鏳r����R�d�Z��@ݻd���V��?ބ���bW �7�]5�r� 6�K�j b<��	I�71͏�@v�@���9um�Oͦ��,u)X&!Q`zJ�-�7�Q�k�)��|X���\�ۊ���������vx�v�0�%�!d�a;����3��Om C�/}�_ܽi[ɲ�J)~�G|��ǭ���/�c��x{�&�	B��K�״p���<��ч(��u<�/q>.�\����� ����鉠���.��$3Ğ���I�l�DYHh~mJ�bgi��ahM�v�U�3_=�G`���U\�A�6���D�|�}7�T��ԬQ�~wY"���L�(|��kH�S������~�VB��y���RH0�����w�B3�� �-)��#7����-�rk+��F���?B�%�3a/������S����fz�_��l��c��ͧ�-�$��m��|X��g�7�8�4��1�־OT&p �xiU�^���ݖ�H�E�QA�]=��w���\�[Ph�[�!���.oE�H����VZ��p�ҹi�1:�!� !���p���©����D�s��sx5w0?�xv���k_8�;�C�nAńJ�]��	L��kl�D~]�*��5/}Q�P��:��v�j]���Z�?�	ys30���g�Zһ�/<�� ��!M�_TnK��X1�}<z�^����~x���]���zB��P���wW��4���GR�+�1�� .ư�I��i����s�+�t5D��
d((����5���d�䯢E�?�al��~~�����hG�}��}��+m�{�lq�G�4Ռ�i��4�:Z�y���˸�Ŗ$�������S��ř�P��G��yu�A�ڿD�6���x��ۀ�-�{�l�nx�
K���A�3v��N��'��Z1��s����#����=��L�����p�ĦtP�׈��b���c���F��潭0��A~t���R�՟O]����<���<��q`������Tp2����^����M�[�!�(��zj����n���˧A�;+����b��uL�����ȵ��`�ĚHt�����3�t��K�8�<���k�]H B����~2͎�ឍ���Z0���[j#b�k��G�~��]_�A�m��j/�Ў����O�{h,�we ������P���.[���w䲣�ytK+����4���xM�L����K�+h���&鄪
��o���n��5����_���qV�7	�	cx���8A��`Y�mӬ
y���o�eZvl<SPfN�I���ț�f�h��u�A�seV��4�
3�?�|*�E'OmѾ޻ߌ
)f�yc&�g,�W�S��M�mϒr���/6�,3�x�f*�'p�n��z����pϰ���(3ꅗR����j�!ϣ�sq��9���H!�g���E`@Aw���ڔ��\8ౄ�q�P�4�&zm[��.0��V�)~]� ��j�P���ڐlg�2.����!Dp�ؠ���eưRջ��ʭR%l��T���5)����,���|3_�6{���](8yk�f}g�W���O���)�+W��B@�q!Ѽm���tC��$�$��E�{�	O��H poe���P���U�IZ*��.�+��W,�:�� Of[ۣ���LS�ﰼ8�[�P)���a��x5%�Y7�=��/�d�����%�i�B!t��3��P *��@0H��e�x^�I�٠K�s �>��I��^.�3���5�z3��¬M�e��j��W/K�b�d�G�ӱ��'�}]���p#;����l��q�:Q��޳�{����}]��uOU6
�q�«`4Ɣ������q0�^Z��;d�"O�/�tȢ`�ED��n�}��o#�OugN9����W�+��39�P�9f���ө����:�$�\p�u]d�b��f��<���bx��Y��v�P��G\�@.0����b{gI���
n�l8��	HG��r��jM]��#�S��x��q��S�nM������58M��9��m�6���}��t͂[�V���֑%�Y4 �?"n�O��1�B	�n��N�6�N�~��L����f��	\g[c+��d�Ƃ�|��9�Ax���k����t@�9"NU��	�r����;�Ҩx��þF���Ra�ס ss8�Cw�pk�:�~���q�(���ȰI�V�d�Ic�$������N�\��������%p�y���G�^����l���o18��@�6��H�m�zu�{X͓Q��l��yl|Bݦ�5)�����푖{ܔՎRK�[s�����V&XgZo{�$W ��,Q�� D�};}}����n]U�r'��0߬ ��+��}�"+��S!�E���.fإz�V���f�p����}(Mw�##���d 68S��צ�4ui5���o {���]��S*ܯ����>Q''[,��'�4y��?��N�+R�%(�h��Jf�l"�^z ����N!L_�qc^I�#D��סB��m'M�����T����LԤ��� A�10�D	���d*�Ơ@nh���!�^��#ق���Z��8쿡+��Y�\���jK��֝ș��kAu�Q�߰ls!��ۊu߈����d2ֹ�g\���+���?���X�&M��߫z/�R$��	-��g�j:�m��9�*�'2>�m<"�@�i��:B�ooǫ��"����}ݯY��I~�b9�q�ʍ��%Ĭ��X���S&y@�l�G�����L�-�|fݞ��$��_t>���,ĭ��8��n�DJ O�F{He��J��%�'�<_�J�*z���}��_�������:�*cǧ����^I�}邌��l��F��	 2�5�?Gq����z���d&�(b~�Oa$��ZWx�(��7���-mk闳r ���h�U�.(x�����9V%ՎBoC��m#H���q��BȎ\8�$_���<r�"z�\pU�?�˿YxV����/�e�ݾ��B��R���5�Ɛ��Jk�iǌD�����O���w�� ?���e�ӳ�]�1�֑��/�z'���{�+���Zb�Dw�M��?�a˦�o�r��V�~�9ׅ�
b��q�9�fala,3��8@�Y,[���Ȣ�&u!O��c\P^���%��w`�9����O�wu�Օ`���lX��\�=>�Wv=5�~��G�)�֪r
��8a�6��j�VK�*��,1����>ׂ�飨]H9̢�G9ހ]n�U���WcCe�@�C�~�а�D������eUsy�j/S�	*?=�nYX����m�i�}�*�Gk�qh;�N��9R��F�Î�
҆�W�����M�,���{���B-�m`�6�h���Qo�xqۏj%�߱�+����^��M�J��N����6h��3� n-H�-)	y#o�2�u�S��ު0vyn�e��
��f!}�+Z���5��ށ��r���>d���)�1=�����;hv8[�t�g�f�����#�k��b")|H�Di����}ۓ�(�(׃�G��Q9��oڴ�O�=�������寵���Z#�,�q��lD���6���˛���˷�����RS�qV(3;O-y��]���͹2�ȵ�w����ZSa~�|9��m��p�=��;j�Y���m�J�:>��8GeJˌp��_��%�p���5��b�`�7A����r\y��c8�r%OO�F&7v��?�,e�z�Y㡿`�jv
��t�黓�}X��^<Sa��ZMdA���Yv}AЮ��m[�z��f4��T�ֹ��%:VdM�$&����ek��I�7�t���y��26Y̨&xҖ���F  ���Zc2����O�\��G=l!.��U4��+#ȐT*ڙk���ۗ�ٲ�tm��v�W������Z��]6��Oj���?�yp-�)6C��u�������MQ$����8��%g�{��Γ�Q��gW�
_^+�����?�r�[�~��9e�����N��/}���d��1�[�L�gr:s�F�OD�f��WM����2gG/�����z開D[x2r2��4���J�!혪I��rf��9E ��hg^���C3��'��Q\�~����!Ӓj�w���9�/bᣔ�7���ҋXDW���$G!�Q�q7N��̋�ԱÈ��YY.��`[�E��KVzؘ���� ]u�}�>��I1"Ҵ(fr�DSY`�,���q����b>�iJZEc���7�S��]�f\[��C��l2����4�N�Ve�2�p4�d�kVGo��a9^a�\pK�uYW��''T֧#-����tZ�>�����ǒћ�	��)��[�D�R@'���E�n�9u���A	bC�M�� �ۚ��1�hQg2���4D��X���n߲��54�)���� ���^I��K^����fA4E#��q�80�di�γW׽�n���Ę>��n4{�3�x%$��2|X*��N6��DTp%/�-�xR�h�Bu��$Q;����ͯ�rD�R+쳙m0FC���R0q������¼��F�n��4�ߝ�c[Ɛ���5��(+��Ru�f�Q)ԒXzx%k5����]�l�e����`wn�XlxVHYEB    2889     400���!�Z)�B�r�o�����q��P��o�6���׃̔���#7�`�!Bk��>�5���_{9Ez7E�J��dFA\�a�A�C�4f֩��p��4XC���{�|�`T�|�g��j~p
�J�z�'濮���*�<�`�9��V��>�ᘢ0�-�8�k3�|R���&��)�Í���w4��9Q��w{I�m�.o�AA1��}=�U(����gVؗ��є,Z;)$�u��Op?x܀ o-�һkCzC��.��հ�Y�x��p��>	(z��w�'��v�`D�����nYk�C'7�b��G7+fa��_:�ɔT�1z��Q-N�
pۙ�*���w��lH,8��qT~���g��j�H��C$����%ɳ��Phj#Y���q�����ҏ���77��ɡA���$i%#:n���%+�~y�u��1
��xg_�X�ı��J��|	�~�5�:N|,��	�&�s_��謯⑏H{�n!�v�puNy�,ߢ��w@G)r�:11m��]P��Vbi�/�%s�J4Ypy����-m���s{�ӞG/���U�D1���aU�:�fzcOp?��f	2�e� %:�?�����F/.�b�`��N��7?FF�%T��o�	H8b
�&�ɻƍ@ݪ�c/�I1�R�m������}=Y�J;�����ڃ��+WQ�d(C'5> ��zx���I<�z�v@^3��d$>Y[�F���4�t�5�8����p�6�jet��D�yӤ� ӭ���k��ծ��!]�o���{�,��D��n���P��݋E����Ԓ-C�98����i��(��zZXP&�w��ʚOHJ��8�А�3� (����?�`���	�����X��@SC�M!�!b�g����}C�U��H�,s���mu���O3����f���"��gIÝT����z�eиt�!~^)	 b�7w��>5w�2l�`&璸Be�燘��ҁ�$p߹Q�1#gӶk'���!�H�����Fnscѽ��5C���N���