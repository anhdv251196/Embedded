XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��9u�V(F��fu#�O�ޮ>�!���^���v%���� ��k��m��G@�Y����RI�k�Ahn�s�Qw@h�:�L=�C���~��6�=ԅ�x|
e���r��ox��$*���u�W����x��X���Nz�2d&V(&��GK�J�V����̀�[1���.(?=�4{0��P���K�����rQ��3@���"��)�ȩ��m-JЄdz�D<���qqz���~�U�t�4�Q�C"���о�����]!��7�|mdO��k-������E ?���6��d��&��Ѫ8�ڱCd�Y��+]�-�<tbE;�R��*���(�U@\n̸����a�űf��Mxl P��%���u�>�m).)[�������ĭ�Coj(��r����X`���)��2y��c�j���C1�%'�
gl�m��K!�uM����o�;�X\wǐ��w�ϥ�iךjD@���Q}���C��F�Yi�t�7�G��.k�.���(>C��s���� Y>>��8LHrm(��GEg(m��`�G����_�&�G�=��}:d1;��G�y���#٪�
�C��tUЅ��[�wi�%ɢr5y.|eYm�ܒ<���%��B���E?��4�7$��uk�S�V閂�f8.�������k+A{���ƫK��ƽQW��%�0\*��L^�c�0�aہ���'e@��z
�b9+3%����� �l�a4e��d-��GT�	BZ���`�3���XlxVHYEB    1491     490t�簃w�>FEl��0Aە��!
c>O_�z^�+	�2c��\�1{��������/̟����M�Fڭ�M�=[��,?= ����d���'1�(���QQ�ݝ�R�9#�f�Az9>�e��Y���\���(<��9ՊwK��j���̉AiBu �zf>R���#����,��.����tvҿ&��O��f�#}�>��°�{���ʐ��}��� 'L����L 꾧�6*X�F��ߐ6uY�Z�G~����ciY��`W��̧
>���.���[ט٪?�_IXo�{��(zq �*K��+V[�t��Q��`��4�X�ӕ�7����A� �b!~�cL��1�?���y��J(�[���{kR
�k�Z���	����k�ch�Fe,z���)���~_/��7ޞ��=h�N�,oG#4!X�36�f��^^�I�N�䗤Õ�^�θ��=�����5ٸ��?4��P��M�	�"ƽ��.A�
�[?ēO鈯r�7	g{D<��S��H�\p$&\�����^ui��)��	�m����N�t\�T��A����HQ�1��wK�Jnr:i��bN��:�=s'	G%�1����e��M؆Dd����d��"�6l>�?4r4�A߈d�}�D��9�
?�1�	䓞)v�f��-�������.B�yݟ{�]9�@7�y*��V�|ha]��۹y"�;��{�V��������@"�~;:��0��3��[�\s�����f�e}p����w40������m]:y޾Aq���x
����l
�΄���6���,���k1��4Wz����7ʓ�����'J�Lǵ�����S)����O��3E}��Lٷ��U��	��>�AӠBr:��(v/j�d����P�h�VZ>�
ߠ���anU��\#�T�#�}$����Ż$�&�CpZ@Z�|�y��.a���I������Q�7�Cbx�-����][�������T��J�C�f4y	�p�^8 %��~�D����r���{�m�;0����	��Ɣ}f��QS����p+GqU���~���"�X���&����<朗��\�AS�)K�}�*��9X`�񠍪_>����7�TV"�*�ڽ�!�F�^�/����EMψ��6 _t��:�U