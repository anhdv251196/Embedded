XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��-f�n�Z竍��U�>#r��^��fr|�6�s�"PG���M	k��~8����ֆ??)�_re��j�z�����&�E�Z�/}!п�d]�	��s��>�T��}��������0�g3u�f~Y��<�_��4`F���}��4L�`1l֤Z`��x�sc|�� 9��y�d߷�ш�b�蜃Ⱦ	�5&�+���WP�ZVb�TP[��Yz��@��C]>P~�ٓ��6R�ܠ;����+�ņ�[>�ӽ�Q�Oj�e&Ga���,�I�}[d1a)g�Ӱvݪ#��^�"F%��UN��!�:�?� AIke���m7�P��QQ����N�qA�7WI$n���l��Z�N�l4FT��H��*�H��չ�R;E����n�r
�� �����C�]Q	^	��������$h�Se&q�{��<KB���Պĩ���h�1ǈTRwaV��٢Rf��4�����dF"�ssz��Y18ˋ�#�LU,��j1����_U8�#dPq�Y��O7�*̃i�m#I|@��%��ZsR `�nW[���?S���XP��v�9�*�ݽN���B�oϦsn��w��-������{�N�	1�;I!BrQ̔�8b՜WSF]���ΰ��	Ey�
Ӹև1Az�9��/V��""]��K���AT�����*��+���4	F�6q��b�g�b��e��@0l�Fl,��������BH�����1���X	��1�_���p �a�\��Q*����4ra�a%�t���XlxVHYEB    5ff1    1040	i��z��	T�����p�P�; �-����sz�*�G�G�<�%=����|���!!�=�Q꜋{��r�V�]o�{�I�X������X�6g<��V(oUD��?���J��J2ʕ81<$���@�j�z`\�J*fVn~��=�(��#�����������`�߳�G���un� ��՗E�
���i���26I܏ᡬ��|�>-^A���YqͲ�G���Y�4�ذp�,��f���/2�NŘzVQ)l%�QI�5���:����V˥�ySeͯ:k���9����o�s�%�`i�M>n��e2NMt)��4^a:R���VWϷ��ٱ@��V�ڟ;�b.�e� �Qĝ7޹�gC&B8��F���;����8j����a�7d����r��Cx{� �4Ǹn�������l�ua9�i�2.�-�e���UPyJ�7��H`�0��F�K��m4աx4��I��y�ĩ�ּ�<~ɞ�5�|����x?�0&x��+-Ir���8}��%���?
��G�;� H�R@˹�na~���3]���P̜�� )� �_�W���H��Ua�Ef6�xo�f2N�d@[T�li��߶�%�Y5��\h_*H��5�وe�r+�	�������݂V��� �*$GH,i�^q�c�W�-���}�.�9m��#;i�l�^{����b=�6}�M񊻟�H�W-ܗQ%�E��ғ�g��}Tݲ���P���޼:<t��_��l�s�������/�:<��\Ri�p����&�nA|�|0�	6-_L����׻��3����rQD��4�dm~���a9q��s�Ή ��<��%�k�2>�Ɋ�HTFE��������ꪞ�e�+@f5�7;�*�ڬ�#0+��&���C�5�'7lK2LC Ɇ��7��P��3*d�a�%94�t�X꬯� b#��yƴɬ���[�� ���<���2��me�.t���dX&��\�Y�6�]��
�i,mg�~(�w,ꮑ�S�7.G���SF�]5�N)��>��������T6Bʧ���݄[���D��î��r��ҢA ����ԟ����G���3��.��U����1nf.���a����ínFŲ7�_W�#O��X�2�J�J�Z�R/���W:t�m��?����7o�"�/���I���
UЮb�ܣ����X���!�E�L"�٭TJ{���z�w%�ͽ���4��_Q�&��q2�K'��@I��.T���C�Ք@�Z��IP�I*�#�wң[@Z
@\@�	,D�U^��h�oij�q���8{5ZJ����<���"	30�:�.}�����lt�@�o�+�D���lO.A;�Od�����]�?�Vl�5�NQ'7^��ZYکXhȩ��%E�{���A ��:��[������A͞]��,kX	hFv�ޞ��
�I'�(���'��y��[p!p�T�nUX=VUO����n3�h�ܞ��u�Cmv��ͦ@�j��u�s��V��ʚ)IT>E+��<�&�+r�mq�̈��;9�'�Ԇ,���Ŷ���>2�/�y?��h���&O�*���N6ł���Ѩ���kh(Gƒ�'��^#d�$�8`���F3�_O|D�`����i��R�D��j,^z9Jd)�Pqd��c� �<ج���~��[9�:	��U�B��B�C[/[�B~��@f�l̯��?�.�۾w�Ņdx�[:��ۂe�-�t)dGszpkÂ=�L�I��Ƅb���n:E�$�X�2�~�)�/�<�PL��D~�5F[9���x}ur����G�[8Q�U�GkSf��;_�{��k�rc0� ?~{/�7�+ C��s8��*5�
�}����3d�v�X8�H}��Ѿ���3�4����|��#���qa-�uz	����k��r�P�aT�?/ �����&�~��h	��"ވ9;��d�li��W������8N�D��p�Q�7 D�xK�wL�w!0�Z�J͂02�`�P�E���L��8�Vzq�x;����oi����2��'�+Qk+�˾_ ��J��W��7F࡬��쉚�6��1ݝ��d��;e�7�7E;��j�	�vi�������s�i6���I��KZ����Zw��"ڧ��B�v�Q�ܐ�2�Ӛ��(�!�k��Rq�#"��@�E����%c�df0Z= �^5���w}J��O��g�斵�O��V=��i�5�(@����xLGBtX�i�E[gz��ϥ%/�".��E��EF���\��n�駺e���Ғ�#V�>ϘKo��X}^R�����'���B���j,�B�����1���|m���k5��P�V�Ɂ��xK`!1q�[#�Kش�"\�2jU���46�����j�1��mG�(C U� �(��8A?�����6B��צ�Íqj��.ӡ�M��.C�þ�ß^�4�LP�a�
⤈�'UX�1�5$M�L:���8%�9�}ս�*n]=���tu��U�y8� �Ʃ럤9�~(���֋���ʄ&P�kܩx����V&���� �={��I�P6��O���f�B�z�����]���I�r�3�J����Fe
��Γ��[�1��]k���ϑ���|�`	��G<�����4cu�� �"��4wN`�AZO�ߜDQz����g�gAyU��&�k�tE�D��^�(98��SW�\fl���8�Bcܽ+�b�).$�6ԡ+z6Q2�H�%�4��c0� � �U9P�3ȅS�Ij�U�C��簠�qv\�5U3�'�V>��Љ=�� <d��{@�$(9w��>��	��>$��D�c��o1͒��a��N�S����fY��B�����:�@�v{]ū��c�U�����4�x�)��
h���K���"��ZbSڴH�'�|bk����R���N ��s�е�n�*n~r��V�A��%{��i���'U�8�����Nߖ���N��B�H1��5SEç+|��y��-h(�3�`ߏ�kp�r�H���{���Íw(������4�^� ����et]S�*�����҈�꛰�yGW`���!��У��_	��h}�V �0%�n��2b���ɓ�*>��L�= �lI���(�Q��oyѡ��b�[^���2	A����8r�?�>��
�1t��u9���G��|G?>��8�T�W������rgz�/$����M���0����Ū��羭���ZȺ��8�W�s����o�V��[�]�j�x���a�`��H/��ԥ@@'	J��:M[��ڄ���p�<�ޚ�$t�+�F��PF/.� ��!q�G�� �����$�^��4�~���G��TD��̦5&�!7�C YB�T�dv������b	���tWgS����"/U�UDPK:�A?7�@�.�,�1p}
V�:E�%+�H������B=7��1KZ���`K&���/�k(9_���>���t��[��Nb�'q���w|	5vv����tUC�����p�hy�5W��˱����+��ܲ=��Oz��6�&'����Tki��Q��,�b��?�WY��9�*�#�}n?��~��n��X5�jELk�G�<��x9K]�� D�C�!Vy�U���+�?�.�_���� �[/���w{�(w�&@9������e
3�8�oH�_N��OC�_%2d�Ã�YTxr+j�~�ǎ�6��wr�pw�|�xz��l� X~?���ȡƕ����nz�I
//>�G�;j�
���NQSǪ�9l��>��-t������t`M% ��(Z�L�PJ�e`w�g���y>1��/��tP�q]9���7�$�I��S{��'�s���JI�Υ��om��`�L�vp|8���ɩy��h��_ݞ�{�r���>-����ݼ�5�P��*w���Pߎ�����2WN����f*�
5�!0��}ɗԣ;'�)
�EQ͊�������@�|4��zXG�j��J�Aڞؽ��y�b+23Ou����aǶ(�٭t��`Z����T1lHiV�ހ��9��#v)��Y_k����.�F%���M��,�s�%hV�>s���. ��ǡ�:��}�t��8�BI