XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���wHqÕF^����h�n�˕�Q���%�d��u$�,�fʾ�{�E��6j>LAم��]8�tJ� �`�A�����iNZ��4���X�]���Ř�Υ��ŝ-k=
���	��ve�����$!#������EMK�za�B��uNB�}l����ԃ9��q���v9�;!�(�n���l��-�.�}��y� �蓝���|Aɣ��MH��B"���z��?z��=��oG�=yb�}�@P��Z�w�m�z�f�X�����I�你�_4(=*Ƒ��2��W��=w*2�l�V�"h�o|sb���Ҵ����m���*f�H�q��X��dYQ��lƛ=^�����|~p�떙������T��q�������.�(�u��"��p� }f��݃�u�=̨�� Hh���	�Z���J�����ӌ`�l�k��(܀߷Y����yo4q,?;H�v�fQ 9�vlz*[���QE���<��Kj����8����V����^�+�C����3��~�(4_:��h��6�V��|aϱl̀:����8d�1F����$nΫo��Rϵ^x
��o�e����b�
Tb$�6��'66,�^m�\�$�AB|�jܕ_��g�;�c��9�S��ӁdM�h"n����ǡ���h[�����|�4�K����p�3E��<U��˂��d�f�I��,� @�TS��r�T�r'z���o�-;�
�d�)�ѥ4N�c����;6���|�����&XlxVHYEB    2d5f     800��q<*򫾛�}P���?�E���y}ߝ���^��-72%v�Y�T�_�����t ��ҝ����M�=e\4*�!��G�F|����"��O���dپ!S�7dh��%�]�ʺ<���|l�㇧�����p>���͑H�n��^ٕ�zJ��p�87�ݦ>��U��V��chᨥ�m�7sB�5&�j��E�E��_�t+��/BS���N6X6R�5��׆k}ߟV��.V\Z����z=�#^�쟎���/H��O{EB�e`�������ѭ�+~��M���W�ʷƧ���	Ռ�|���������&:Zl�'�}PS#�j*��F.��"�;<?�#y��(��i��u����u�a�$fsd�Nt/bi�c��ה�1��F���b�'l�ݟv(��6Q:WG���CbMjT@g|4���Zе'�nyR���n�j��U��*Dx�1bBy\w��]�H�z Տ���y5�F�8�	ʷ��Yʻzx����|�aE���˿��>9#n+��x�,v��x[%���Q�Y:XBe�WZfof�Zk?� ƻ�o0�\�^��tT��]��o�>�U�E��P��2�S���X��RME�R��E�E�(�� F�0U�U��l�b�Anġu��>���`�2�mB�`�>��z,c���k���bq����(��˿qܬ+r^!����q�p]�=$��'ڄ*��Ӂ3r>g�i;�� ��F���|�i	#џt��b5)�Ĝ	���k�}g]�ǟ�3�D���b�5[q�jdhiVGFg�M%����hۋ����݊��|(�M�b���E!�J�Oݼ�1�Rj�yh�H�om�MpW'v����!sBN�Ƣ���E/l�=���}g:/���U�U�����>���Edɺ�׼��y�2ĵ��
x�ڢ-mdjE(쳹��̥�z0���Px���Y�?�y�I=�+��;�}�^�_��O�����/_�QKIX
�����/��-�I�-�% .m�=��4i�~Wt
�m�=lm�K.��>�c�h���7�b<���q�$��yK�~h��"���PX�?�U4��<i"�pA!�(�"��%Eء!�IT��a \~e�>�������]L���=���8)�6N<w��e���X��1{�`/ 32l�oRt�iyW�b�f]i^>,ޥ���F��Έ3͸����*;��k+��N������FO���';/ok)�v�[͋�k�M�a���h��0fK ;%����	���ڵh��pņ_�'�깔g���x�i�A�eI(�wg-o�*�Q�TJ��7� ��e��>᝚q�;��<�!J>�$�i��V}DFL z0�0;ǲ-�ܚ�{e�?V��'݋�ܫRY�=�PQ#�e&>Y�)��4k&��0��ˏQ�[��6H����I��d"x���Z��\E�lH� %�3	����r^�py��a��[$;�JZ� �4��U�ޢ�&]�'G���^ƀ�qx�X�X�{��~���X'��<z�j է�E]��@�����+Ѳ��>�,V �.�i3/g��;��'�v�בB�<�/i��1��˖�2�NP]`�w�E��?(tb�ɮh��BY����C��f3U����wh����@K�X�������ʹ�(�a�D5�Q����ԓ�xX�Q8��s]�f�d�w�U!�U���/��vj�-ǘ��P��QP?���`h��I��}����A��9id��[���N�3���k��΃R���Gf�儐q/����R���+��k����0^��"C9��%;%����Ug]��=������:OQ��j��-mT�y�c~�!�~�!p����b\�^�9Wr�'X�s�rJ4������\ߗ'��f�}�@Ҋ9�=�I�|$7�ؗR1��D��Kpt��7]l18=ڙ ������!��re�<�.q~�����vދ ��Pn�vz0Θ��ŵ�E(d�>[��=�9�!�<�y���Ni��#�jS�|�<�0�&>),i��*AM