XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��{h	��~�F_��X�U�k�A岠nw<MdM�߉��X	V,Ī��<����|�o��`W���)�s�=v�H�?�Ɩr;�joc/S�ww�̭��-��!�>���)h��:��ܗc���+���u++}x�O2���J���C�������1'�n!S$mo�M݄u�Xд�I��όF�L��{��_�5�
 ��Rd�4�3@n�c�|�Qt��i�/��,��c�zʷ�������: Q_ ڴ����Si�1~�]�5i�F�����F�	�i'5���7qDzkC��c�H.QC����kG�E����(jux[��*"7� ��+Y ~��=aJ�������r���P<�y��fѰ���k}�P�̿�������/���gV�wxy'i���`�o���D����h���'��HB�$�'�ޞL:�N�,$w�\:��.h�7�q��\ee��q��s��m�sq�.������a��	�7v���?Y)�d��F�	���	b��*'h�'@�n�H->�n�~\���TCF=�
S��+�R/����>3
мR�9aLI�a��۪+�a�%�7ݼ�"Ѹ���G���@"�W��y:�ʴ����P{�U�̥%l�!�
��T��l����1&���כ�V��[�+wV6$������o��k���j�Ȋ�Eo|$n�z��zâ5��'.j�O.j[X@ˈ䉳R�YB�u;�R�0�5�0䧚Y�Q�4ex���#��8d2����`<TODb?Ā_�7XlxVHYEB    3a1c     d40bK�P��"L�?_i�k=�{L�\)��Û�jZ�น�r:�U����r�a����<�����*���u�)F���k	,��)�@�U�G��-�a���m�@�8���?�8�0����n[�uu�W���ū�Z�C|e�	����ii���8�Ne>SG���3:/XZh��(�����0�Z��G�ybA3���rRn��c���͵P��a�RCz�x�.��p�!|��t�0�K@��-��а�/���Bq��B�w�<�1B�ܝKI�yQ�,��ӣ����~?~1����)��,vhU�3aH�}�F�u��݀D����#S�ɾJH��M�.�g�ա�{"��b�X��&T�(�fon�T��%�&Y���`�օj�uI��u[nNX����O��8���c��9Ɖ?�|��J�K]#�޸	����u�L�3������7^����>���ܷ^Hػ�3�z�� ���OQ%�\�I'�y����~����s�|�4,���#@��k��׵r���h��$��O���E������[�u �a�=F��ܮ���̎iuC����CQi�����ޢ��݊YV'ڭ��{��@�b@��Q9�^�Q����� ��O�|]�A���%3����R�/nr���x7���:�3���b���Y7��ؐ�ף���恙����(���\b�����}�Y��F]��<��Xb��>=Sk��=?�[�sǓ������NY�2�A�ԥ���N|v�}E��G��T��q;GeR�
��v,�0C���sT~�[�n*������@i#��ҙ�|t����!\q��?��#�e�@2[͞�`J!w�".�8F�}8~��G�*����69�37�3#�|=��!Ty���Q���<���Y��3�2�(��}�pƽd�Z�@)�� ]`W�nV5&��uS�z�+'�B�߿�6��m*�w�dj�`�h77�Xp��l���>a�-�[�Ju�.�� _ems!�H�<G4���5s��� �*��t�w�M��m&X|���BV=��wIY�����`�v�?ȿ{`��U�P{6ȕO�^yU��<�UP9����z����.�:����)v���+�e��l���I!U�e�d���A��Rݏy���#XJk �H�c��w�������(�U�*��lV�z�n�IF�Q����k&�_1�B;���S�7^ɕP/��G����q]�RaR�FI�����%1�!�l����S�	��jT7HCf��;�~����e�/)��d��.:y�U�# ���MZz^
3���\є��F
�.>a��7���X�Q�G�D�d�HR������Ce1�v��͊��Z�Ļ5ȶXH�=~# (o�����Ln�h� ���M�%a]�[(��׺�Ey�t����n����j9`l�|����G/�VŁv }�B� EB�����4G�.|AM�_��58V�$2��,��}�բ������s���q&��^�)�b��V2��.����u~ʳ6��b�3 ��cB����V��-�b䛛��S�aT�UF�|�E�Nf���M�(�2��H�%��"�!���3�@�"^�J:��k���*4YQ~ ϳ6�4d����p�5�6��Y���SmĨ�S��A���c��l[]Sf��c�B��yh�=��6���"Q�{'�|�q#������kMʙ}��&����p@��X��-c�jA�
G��0�����]�)΃�ID����8D *�6��5�����mW|��%=�rb�b��G,�$�9�}<	>��L�f�-�����k���\?,�g��*�P�k��Q�\�.�Ɛ����A�l`d�Y�O��t�I�r<G~�f�zv��UW�
<Z�e�/:&;u��9��p�%ӳ=G ����	�F����c�x��g�����_�h��գ�"נo*ɵK�[�L譔���t=����Ql(3m�~ǳ�iVK�y��뱈�Rđ���c�>��u���#uj��o�ڳ�!�)v����d�e�V�z�ܛ*J(�j��Rx1y�#Ս��z�����#jFRA h	����*�	���3Q�r"�-�����|��NO=�P�J9����q��@,{�_ǝX��94w2�k����Vf�Ҍ�+}�jg���NK;灇
oLXn�er~&<�
f|m���%�罆݃#�@�z��x��x�T`��yǹz��Ů��Mq�AS��TMM�0�K�ѫؘ��>M��zh��/_�\�8`K8����i��)�2ʙ�ɬ�$�%�}ٱ�>�f��G�N�b��ѣ$��@T��_v	��Fzt���5&��4�����~�̄�MC��8���2I��	��N?��f��&CZQ�0,��*��q��9��;Մ_�{�HQ\�����
w	���T¶<y:��E�[#�2��}jL�D� �3O�2��6��0� v�\B}�����/S�h'l�h��*��V6�u��	�`M���M_�Z��&��Z�iF�8LN'�/$�r^�%EEof�ǌ���'��~��9�� ��=u~ָ���1�Ͼ�g�G*��~h?�j�&Y�ɚ!��4&F��hkp�5��M����v���`)�9���ʃ���g�p�:���`��3��@s�����Cu�;k45D-Ʊ�e{e�Qe�"��	*2��k�K�N��s�+�e$Wd�E��G���K`���sdM*g���w�I��ή8�k�I5^_�����Y�n��r���{�GU?�pb�VU�ܢ��mޅE�n�"�����Ҭ�?�(;��7�F�G���!=(rĬ�S�|1F�j z�k�A�l�*��	��ѫ)�>�����2A�&W�~�����0���<	��33��8�G��!�	�ZLM�݈��j��e���Χ_���#av�B����QZ����+�|&Eφ�3Nꈾ�l��C��)]w2I͂�C�8!��N�c�FR�V�����n*�f��������1z)�X��ӟ�|1:��0)��m�*�g�y�U���Ѱ��d��S~<��H(d?;��$��S�23�%n����L�'/]2���Y��.�����1�juT�[c�綋安�����[�Ak�q�ȵ��?�>`�7��]f��>��m���H����P
��-s��Ԡԓ�2�U�86�s�m z�j����V,&i�m?�u�'��n�A!N����"q���b1��$�*��C� ����[���1�������C'Z^0���ECNq06��mU;���`��K\O����coYPT?�v�LЎ��M�ʑ��cnt�?3���/��!͛Xa)���3�P�p������Pq���