XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���f��:r6��������&���	���~�6W�-����-5)���B���zQ�O�n��h�Y��$���W�YT��<�`��(�p���%F�C�i���;��Ⱦ�j��a����4���z��,3s�1
q�(B������-�l���$�'H9[�����1c��s�2S[�0oE_\v���^���ؗ0�#!�xtP,+�����KN�O����Y�jaIb�=��4���t��U͚�N��a;�c�`fW;���z'
�R>����M��
v �a��c�FM<�����{֟�q0ʫ�����y�<(�c����@�<@�/�%
w'�O�T��A�b���o������ط����V)�RU�	Ix�R�-]0rF��y��D91 G��1^
�F'�f:�;�<,0�+�!��%���6'=h�[�2�$�7��V!��E��7�V��>�9y& Q��.��L6�����H�zEMH��5�3 9�/x��I_��VNi;�N(��N��74��q�t��^�,n?M���Bd����ϳ�
dɉ6t4ʨ�%/rTW�^ZRd�:���h�L�ê8ĐшP�f�����y�H�K5�"^�*$! ��V��Z�E&5���._&G��C~$�_@���s��
��X��t�Sճ��*
�����y\��G>�*Md�`���z�JY>=�TE�����9}Ĕ>Ң���q�I�r��QB�i߯���F����RS!")��wUok.�/X+"�!�+p����XlxVHYEB    1cf8     790K`�t�5�����PM7�'�Z��؞���%�^d51]�e���	ڰZ���k}���6��Wq<evLC����,��q�}���0��t��>�Kih��p�.���꜃���;�Ry~���>J����b�SA����!�jvn�1T��0x��s�Qe���G~ �������[�u�{iN�@�^��$}p��BN��ޟ�ESm�U{/�z#D
ݫ�Vo��s{bma� �X�9��j��ٽ���\��C�(@��ʟ]<q��h���:��7T�-���.�A_:�O��Û'�.�9�m�z�NYg���0����=��wJ�v��gyuR̬����Yq^0)&��&n�v����E.*�ti	� �.���c���3�=�� P���K�x2�(0�Ƚ�,u�T婭�o'�(����Raڻ��tp�j6��PFG6Ap	y����*��#Ċ<=�jQ��%���¬?��.�@؍�4X��z� f�Kgr���L}u��7����|&�dJ���D�U�b!�-���>��l�R�zV�:�[У���[��n�]WO	�p&�ViZ"^ˍi(�3��_�r��31h�0;��iO��"�����ѩ����uq.���r?�//oW������1P�J&�F�K7��>�NT�k_5�a��P�&:3����d��u�J>�u���U� '�Q�-ů#�����H�B�>f/˛��5�H���������z`�Ų��o:���hq*! `�U����Y�d@�X��|~��Ӄ;#�8ta]�@��|�@��$���d
��r��]����da�m��]<�/DI����0u,�����(d�`�k$��L�r��������^�6^��[ѵ���	���Q	����<�7!H([��cC�Rx9O���.!�s���F�V��˭@)0q�4CP�a��i���)V�߫4:P�<���5yn�B��SE!���-f��x�O��E��&/͆} �=/|ֺc|A��W1/��B0�<SӸ��"v��wD�ֻ;��j��{�����ð�mJ��1:�ؙ�2�!J��p�l�^�
v�����h].�hq�ke6�7�1��G�wr��VQE����5K�^4(�}�t�Ju@ޒuj9:^�KJ�0O%��P��� �qoeVDNs}m<�6�p�����&�%<9� M|��Ŷ��'�</��ǡYܦ��U��&P��nۿ� �A���uh���n��$<����D4ȴ��|�C&i0�q�T ���B��q &��Q�j����i$]�	j!�7rD��W3��Z��)#� )��o��bఛ
��<��w�����?\q_�2c�����J?�:PdB��o�E��2LW��_8|�D���R��3��G"�.m9-v�q�Uz�{�dKn���߱qT"2j":����:j
+�'	�s�3���]N6���;L�b��rxonc�������KF0X`���F�y�طuY���C��$̖.�r��[*�$��l5&���Nd�Ii��Z|�T�+�jZ��D�MR���R��n���F��h9:�s�Uk��eZCIe ���/�����`��i�b���ʉ�j H!�d2��9�9�w_B�u���`�e�d�.LG�s.�i�ў5�n�6�
 ��6hݣ@�U�qڑ���@@�0$�� 9��t�aC�U��#�CY��Y�L5l_���+��jk���d���f�l.ߗ*�'��2����u�aA�I+�3[�{7e��s�z3O�r�#����t�Ms&�Rt�Ӿ
���2n�r�nAʙy� Ghd����<�S]繗�^\�>Z��$����(º#P��P�i�]��o��u)h:kb+�'�}#�o�ual���ݸ]��fWf]"^e�?�B�Hz���-NȻ��~֛��{�!Ց����ˋ�f�?�m�ˢI��