XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���a2�4sHq�9$A��\,8�*�u\u���l`{V��I�� u���u��ḕ'OC��xq�#3r��%+�!���of%Sf�?� ���ր9�{�6����RZot�pU�A�aHK��U�{��]���9E�o�һ��D�F7���R�C��*hW�X\~����+�A*���S��Ci�JC�u��q$y�Eka#A�h{�n��n��-���G�imw��f�y�Nʨ7<�M���s���b�x����]����V2K�(W�Z����.�Ya��׆Gb��r�L���G@常S�ä���^�'�fۻ%ё��J|/ﾆ��b�:��t1k�l:�^;��wq�p.D́4��9/���j�pgQ��Y����%פy#\������#���L˰���O��D�.\Ɋc�?ɺ/.�@���t����D�%�)��l6�j-�脎ݡ>[�\�x�P�+@Q��n��d��8UA�0�fF�_�0˵e:W����Y�9�@�M�x&j4��� ⵶F)�l��_�DԼ���u�T��o�'2�2����]#�E���d�� �U�c�ӊ����%XY�]*��rd�׋�	�8��'�4����8��4��r�LM��R�d�$ ��J��v�~yT���ͬ�߼}�/b3:ڨ�D����aY��`E-O���z�C3<�G�G�q��������h����%90�,=�������̮2�T4Is"׮,�����pä������D֌Կn�E�U�Z�[ܩ�P0Ը.��q�XlxVHYEB     705     250z���=Y_�L�6����Ņ��9�Z�z�K�BѶ�އi#w�6W�D�<ۙ{u�������Q{�cA^���M!$����]�o�z$��R��؆d搈��6ڹ�.�*/��7�<g)t�b~|V� 0�IB;Q���p�^	^��;����O��N�
w�J%S}�E�h�#�X�Xh������r(� ��!��/�P��S���P2�8�o���f�9� �?	�������s������qs�Y��A��x�e�v�8���I�ߓtĄ�F�|�:+��3�Vs��	x�u&_��(�Ԧ4�rNidc�wv�n���BC�(�ˋ�NpЎw�%�k3�cf|��3����΍mW�o�
X�F��)�f�
��;6@�F=��e3M�t��S��\�]��)�%rռ�J���w��!E�S`lF5D�!�F�*���skj�@�7F���1�)��[�"�V�W�����J֖�H?wfӗ��ԙ:f
���?��\~��0Ǽ�+�嘅��6!�9.5�h�4V
YG<յI��q���ٌ�r�+j�/�EG{P�ص�ڕ7���.����`D}�Yd*c�gB