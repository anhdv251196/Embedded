XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��[H'�1�/^�W ���w�^D�'�J��!�-eH��#)���ah�p=�t��ֆq��}Ӧ��i{��+��'U�/��Ka[����ǚ3���7������9(���^�X�&��8640�L"���~#`��h��Ʀ�-_�H�A{.Y�H�L��J���������U"�r�}=2ҍ�;`j��%cr��`��
�\Co��Ru*�S��ۙ�<cd�����D���aS�?E�Ud&]W�f>�̲�B`�䃡rӬ��Z��.��� `��$mi�"0q�'�y�I4`c��	�VbS-M���!���5��W��1����`I/�H��I���FxT[����ٱ-��&���h�g�ǅ���P�Y1��c��[,�p���DO���_~œZ>��<£����t�����Z����I��k����7+�\�ی�D�Sźb��1F{�s��� �ю<��Ϗ������ߛ�a�_���n�;:r�(
A,���!%{_�́tc[9��2�2̬���8/fb?�䰾��	{qЯ,{��$;��B{n�B2��C��������^>�w��G2��6?\�0�qu�f�%+�����Oeg��������Rd(���*�D�S,8�I�&EY6�âȇ����=���}�����M��p?&�4���p����H�V�9��	�gZы�o�f����
F�%w'ߏ�w����?���Ŋ/����	� (b�]>iAP_,��y�߉J)r"��ߠ���LlXlXlxVHYEB     7e5     330��
�{�x/��|s��ƣz�H!doǂU_Sd���;��צ��;���+�I0h�M�ф1׮g�=8�Kr�b�{�M��k�0�8����R'	q!���]����jc$��("F ���W.��!e	�����q�t���Y�{��/E\�I���C��N>S0�wYAz!à�<R
���?��|��\��G�@I&ew�d�I�3���7��ଳ��ss�&���}W��<	�!P��e!�8�+a�ß�T�@�g�q�L��Lx1���ѭ���ܠ����"mso�#��n���* �����9;�O�q��� ^S`�p�L����oL�k�pi�-}´*����X1�A��z;Z��1�����yҭ��&���i�;ā��$L�5$o�a������՟:�^RDp�B�lzX��/��(�Ya�+m�)�Sh���5��k��qe.�M��|(�����z��IQX�_�KQ�q�i��s�
�=�_�
A]�!jV�
�x7�R��Ot�	y�P�s����0#�%]
�'�]�ݙ�0H�H�#݌L�ɍ/�#���]\���(K��X�a1�T���-�{�V��֓J(8�|<�����Ke�7�8��%5~�W[�m�����`҄a̭"�.9�.GbN9RA}���_/�!G�@X�J�x�qh�Q0��h3 D|PFc͹��u(���Ru��OM��v/�W/���r��8k[�R�}7��{�Ѩ�&m��h����E�h��ODvV�n6HO%>��k)Ў�}��b�	;}���#��r�4H	��FFr��}���Pr�