XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���P[�͚������yBM2;ʘsjFXߛ0�K�S�s���b5�J�5�J|� ���1`��E�9sw�՗E��
�w��z�O�K���A%*��|�*b�d4��
9��~�K�~�~叾�6�\�<G��@�9B�@Z	�qP�`��7�@V���E��P�����c{_؍�M/�-�%v�8� <��o��)���S4�Y�E���!����c�M�����A����_fp�&4@WQ��b��a�\��'�w�Fw)�B�C�B{ʸn1+�N�����SZk��,�����˧A}�TzJ�D.���[&�9}�J,^���~�H��1A�]����J�CT�-��kcI����-v��O�xk�H'�Ę�2�V���X�B��У-<���|���"����0(�
n��|"����z4���3��5]L�N���ٽ����=�dο�L`���]���ܒD�l�����R�<���'�`������r��{��l��p<�"XO�(�Gp,��9�G���@����Ԝ��d�#���9�A�R�n��4�Ǳ&�0�����0��p�~��?��!�^_D>3c�E⇂�d�Wl��%�2!��о�Q4�LjT���tn��G�)Һx���������n�V�gSô��U�d�m��b� q8B|�����j�F���լ�f�Q%�A/���8R�^�~�}�#f�I��vd�E��Iwڪ�d���Y>�J�C)1��\Hd��i���3����"��
��4ۯ��XlxVHYEB     9e2     330��/2�+"kp�~�$\Ti7�ٰ�VH7����� ćڔ�x�ˋ���Udg?n.�Z�
[��i���`)���v[j�T�.����Y���<�H�"w���7i`Y��<�<=�V�Dd��y)����h��rVDe��%,R1X$٣��.�.�]KJ��]���<�]~ŅDa�ϊ�b���v+�^��o^������RQn��U�|���|��ף7�#a�/Gѯ\�}H��
=��ݡ"ꗅpy�]�LbN���E*lfd��H}ԃ=g���A?��p�~d���ۈۭ��V�T{]j�W�o�[p.�e� ��$�N�#�ؠ�Xgv%)����!FKk
'Eq��FbH,�m'���+��zˌtd��Yp�ف}o�A-(�:B"x����M�|�j���Cj�9����O+$e��5�s 5Y)p�l 	��t����ڝj�� m��;�tw�-[��Ě��RIO7�",Q��3}|W#������.ڢF����B�c��>aۧ؛K�dy��^������h�I�Z�𑯤���kՎ-��I��� �����#M̹�$�yT��n���/h;�Ua��D.1�@//B����kO��`�sU �����^u�ʘ���w�30W���˧�x�w�^�Y��,�G��VውV�m!��9q�=���\G�i����fv�����W$H{�1�K�p)�0��U g`v*C�[(=K@@����3�E�-�c}���:[J��^�C�F��+�����f�^��I�'ʀAz^���^�I��G%�9�Nl����&h*O�� �>�Yw\d��