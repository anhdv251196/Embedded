XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���ߘ�"c�C�	9�?X-U�6�k-���D��9rew��:P���&[K�>����u�#v%�yߨZo!t^�|�h)�M^����F�׻�5QKeR���l�Q�`��t͒[V��9�I�ړ�`E���
�9��y:�Q��C�o��vE��nXvQ�]����@���[�O_�Ъ�eA"[������]Ȍ"W?%���_����� �B'���h��Hw^T���,T���ҿ�ݦ����]�}����a�h��!v�0@��%�3-���u��'�[�M�p�o�V�v
���~jq\�-�H��/�(�&�����؝v&�����VE�����W���Ρ/=�x{��`��:[��CL�D �+��Td��B{9x�o���K'�������`)�/(*��+߆�pՉq��d���׬���@|�s�c��_K�b(Ǖ�)W���Q��OD��C�Z\�x�To;�
x�isc�#S[>՞�68�â�%76�
�upsq�7~���[����
�?D��Mt7���v�\*00m}0}�u�,;�0�9���\#�
�����8�(m3͐#3����	��k��v�!��%����sfe��|�p_�QOK�~����*�au�_��Ύ��'��(��5W*,{��4r��P#���}Ө�-)��ˍ���d���=V��rVn�y@����q1_$�������5�X� L�X��� |�~�w3�:���l��DA�ω�({U�ԫ*�q�`<�i��,�H���XlxVHYEB    fa00    1a50�7RS{K��(��túĤ��i5��(�dֆ}� n�i���Y
��quЧj��k;�����-�+�.bQW��9�]�~=��Y0����,����n�A�z�¦(Sۉl����KW���R�ׯ��^���b^�o�V��R�/�6�;ZI%R����t���9�y]ɦ7�I�#�T�9�r���7��w,�?[KM��Įy��Y ��L��	
���ZYEm�2+�֣��`��b��[���f�9
���!ΛN3d�Vf�[��5w�~=m�͍1Z�_ʁ���7?#1*	�-���v1�����m�,@��2��4�wz���."��x
5P�g��<T(,��5��f��������>�퐬Z!@ԦУIi>�%�#� F�H18Ơ��f�3��2\Uǣ�KB���F볛	�]ټο��w���<�xc����Ľ+�Xp_ }�]E�J�^�p�s�]���70��ǿ������M]������W|	��y��ex���Ô3mO��i�᾵.�񠜏���)\�kH��d��c���R/=}�p�
{�Q.lʹ�p�8;}g�,�ڦ/V�Zs�ޭ�.B�0S�a���\mSA��dT�i�a�L�n_(�Xe3����#c4*� �@`�-��;�V��K�$�wWu�j�D�]��Q]�خH+������_��X���RgJ�ݶ�Y	֘�F��]�|�n#�	O�T.��b�����z�"�w��|�_<�Xd.S���Y���T�n��n挪��.���X1_�H�����FM� �e�����"q���.<�hΤG���)��]O������[���r��e����+��,h?����&�k���h���G�╃)k2���M3�?��}���.������_BhD׀C�#��/�n9|�� �L&��f�p:�]L<M�ѓF��B�>4��UDL6���4UE{1������4�V�}�&���t�Wա�i��wdi�F �o/� P$��8��i�Dm��߽�j�-)��rI�V�xնX���t"�'����jv�A��J_��b�j��p�k�+q�	����o�q��]c's���4j���D�P�
���a�1f=��So�6��90�fτ��S�w�ȓS�*�4��Ԩ��:���4�
�4aG�3����:�7rx�S՘zB������F������~����������H�2�����������Q�ڟXFxx(�a��/�a��0>7�r-אj��� �ᶧT��G�"���Pו�xLώ�=*V����-�vt� n���!�]�/+iu��R]�	�h�Sݪ-�8B�&	�)�2�MW"�-���2H�E�=69e��LBy!�Ν8q���ݪY�SU��f�r��@s	�V���5�	O�/P��, Ϻn<C{2s����d,���Qf3�}�=��'TD�s�L�##}`���)Ez�D����.Ut�@k�F��ŗ�Ja�{	T��A�����"8;$RF0l�2�'��oB�/�I�A�����c��g��T$�g�L�q*r�Ð�^އ8r)S�F�F�^Th9۰ȸ�bH���-��wq�
�hK� ﰺK��s�yZ��m�p���Șz��/���'����`v��^� �ߣ'nEgM\RUU��k�:昑Y�����u�SZL1�s@�n�쮣�-�JlZ|Vi�UH�W������/|�C��Lf�F��'-���xW��l�3b9�����K�_�����:���X�vZ�U�a����,�C6�ڷ��@�0pBxp�����QeL�N<�鑮~Q��$��])�h<|�����\�yw�ǿv��J����h�d���m�߁�����S�X�|�iB���c���
�����VW1������{�g�e�
�H��,�A�(��0l! �����A�_���7��0�׮�`�5�e�*��M6��.@��-����H����-"E���d��3�����N03&ħ�6A�"�8�P��.tU�M�:�����h�ԫ,����.DU�"eu��j�X]�n�=��u{����Q���T�f��<؎�o�K  ��Ӹ���{��/K�������\K��J���i�z(�4�I����'�u[���O���-3wľ�u$E@{�Em�m�?=	Q��7�oJ��5b�&�&�sZ��h�W�a��_���nhjp�~�$`�a̱ڽ1��YT͌i�tβ ���AuM�{�2�-��qj&��?����M5pr��:4���b� 9�k�S�Y[���/���Ksv��O�U��!�Ð�B+=JB.ĳU�m��Q�����<�m�¨��t_��(�Zf��N�_D&�cp��ಉSJqW����v���S�xm��r[�J_Ň]b��;�����ͳ�z�9Ϸ�Ko����!�	_�'}�`�'X:��bp��X��ݩq���q�ڳ�����5�)@uåT<`��FyNbI)�2��U^� UN;��x-4H����{�@_P��ŗX�D�Z���D��M����Wß�T���5��U�<j��^%�B>sM�A��tr����o�j��Q�0�4=[f1���@�ő0#1,�b�л� �P��j�zx�y]��{���B/��aL��2���[�z�
2�����j�����.K��viN���X��H�}s��雄)i���c4�a<�O��B�S�]���wd���p�Y%���)���+$w<�aI��>]����0��u�Cc6L��؃*)����1��%2��xȟe �
ݭ��oxY���g> ��kǫ2�!zr�1Rc2�#�d����1n�TD)m[�y��L�ē�g.�\��j�CF�OĽ��>�cBi|��K��-(�f��-)�um�:��p��)SU�>[����O�ƱTu5/[3<�䌱U=�D�����@��s����e���+��j�ɀ(��W
��zS�Q�w�N��#�<d�C���U���3�/��d�B���
�#Af���?�N�a]I�R���a�<�'H�����6�������d�1��<�D�b?0��#R��n�k�����M5o�p�t)�|K��"qcj�E�rS�o���VA�%6�fU�%QR��=o���I���Ϭ¯�ӈ��s$�ᱪ��1.|H$�B{���H��U������$�ܦ�i�6�C�5;s��ӧ�6�)���2�f���cQ�N��@ͯ[�>7m� �¯�3�e_�<?���`S�KB�$a�:���Γ���}&�j��,���T�[�-�&�Y� �/�����N<�y�
a�8C���?�0�'hY��O(>�;�V�����|����2kw��@���M���$��V7x��7��� �-�wF�n��'�vy�*ܾ��3��)_{+���lQ>j�c�[�����.S��e޸**^hQ7�S ��"S����-�`X�(����#�NN���o��[�ƒ���<_|�����mN����k����ϭ�[��J�.j�]T?���vFI��9U���D�lzM3
�S���,]���������������S�i��G�_g��W��{=�T�j(��/���~�~ ����m�k���*���d]^f���Z��˗{�>����D���k����,�-p����e5�`l�5�zm2%�v��gx��GT�Y���M����y�1�Y����Ib^6-�.�!ԡ�´éG͕�֠OU��Bl�W�(76� ��E���;y�&�p��b왏�z� &㭡P�c��C͈C����wY��x�OQ�6��HS���"�\py�w�������<I2!˨�R���N#+$���������v���s?�a�&��8��u��YBy�rf����B��?����qY�P���9���2M�[7�;AM�4��R���@7�v�u��r��;��.�WX�tK�Ġ�Ԟ�2c�#e
[+#�����H<Ǒ��)�>2�i��FW�WB�V�����k�t��:6�i����j ���5ǽpC@r��m7U#*Q#��e��<�)�ap�M؀�ׄt�0|�U�!F���~U̷A�*���B�%}ޘ������O$uRH�`5��R�Γe��/��,m�,sႲ�����V{κ�?��Ȳ�I5Z/��t/��Iugİ�RP�̞qCB-5j ��".Cx�NO~2��
�e�2g��t�5c)(c��1)�!����dIl����-l[4+#������m�� �h�ǀ1�8��؎A�l�U��l����������d)��p�a��zH��3����~�R.s.��Ю5�~/����z��XC�K"�ϲ_�cA��ה+��?�귍�6ӻ�A�B�SM�ٝ/.^�Xx#q�볚 M�9���~��I�N�������\�nӄlj
AX�i}�hm�t��g�+��m�*'.����t����R�4����K���d8����j15���k����^Ma�
h1�|�*�����MY��%"��eiэ���o�O�d�����H�J��|�׿�Ӫ�x"W�46l���]J�;��*Tf�lE���)��6�`�52�����.(�ȢdϦ��7��@!tB�-��#�H��M��GW��I��-�Nl�9?�k�7T���ӽ�W�7�j��ru��L.�,n?���2V�9����i���
����]�-��ډ�aSJ�tF�"g���N|y)��!yr3U���љCa�H���EM�$��q�x<p�n$]��T�u4	��mBQo�a��$��)}��V4�hK�Fnfᇶ;�g	�@���ۣI�|�|*�9���ڷ�t>�3�&�D`@����#*���^{%V(��0� $��9�9�8���W��ҍ��U��͌n8�yX���JH�6�߃<_�`�Mg�ְ��A2�͹��檀�u� w�]�2��,�3v��-�*�?Ƅjs>:T���B� ���&`w�6s�H%/��#9����I���͇���`��]�O	~���|��&K}�mzbob4�g1�ǥ��P_�_ؒ�c�KM��޿�+v�B�{ �¼�Z�ɢ���Q�9V�O�?����z���m���,�\D�v,]7���/[�V3���*pMg��\#�2�����{A�T� ����hw�j(!4��g��. �(�||_T�/I-�!|���7Gk�U35��`?m�K�@nM¤�Jr��b������Y&y�G�_2�p�C躮f���4͖S���o� R�z�nK�U�c�ɤ�K��Ϙ�����"��䯹�-bKP)v� ó�F��S!K4O�(�Ξ�:�lk	�Ǫ��*j䰟l2���-�
�,;�{�?�v�����֡x�Bw��z��T_�ĳ�SЃk�k���a�v����}ZA߄�(@Ķ�V��}o���ZT�P���G���ԝ��'��o��+�?�tz��:\<���?�<�%��zŹ�H�$G��
d`.j�-j�-
%�#lf4.���`S �ཾ�R�BM�{Nn������>��e�j������Ѣֹ�w"�S�����{���`m��A��|�8��n��)�S�Y}��E�INz���s)F4���(���7��Y~>�;�� �M^+o��n�;���'�U�X��W��B)L35(И�VP¸���#�ڌ��%vh�3c-v~:% 	6R�p^	MM�?�FR���i-��&uN,�t&���������w�S`��pK�4��K�Uh����w�AjY��d�� n)9�B�G����2V��ﺴ�;�d��!����W_^�h~op��v����x3g+�,~��ޙv��٢��Q�k�X�!���E����)�e	�q�{o}�N�Dya�P��:l񩐟�����vS����Ϸ��kTʸ\v�3���Z7��(�4~L[��{hmt=b\���,�	������)���X\���*��?��:8��A�/5[U�$�~�x��q��hzų�8��=n!��N+��0����m�#�e�#LD��k�>-YZ]W�srFv#S&:(��2�(�7��������rb�Ӆ�@C�p�S��ٻK'1%?2��$��솥K@1�y1d�R���� ~J���q��:�1���JD,Aױ�Yg��y?E˺���гEW/=�E�n��Ivd��0�x������R��6��5IO�x{�(88s[ �C��gp�\H���Z~okY���[E2E#lk}��"U��>�؛�z�|�B��2��&o�������i����I����3�Ou��sj>&>h�
�ȼ�`�E�ň{�/^f3�5���}��5��_���x�n�3w�~�M�>(�#���,�ZQGI=�\�Lߥ'��yf����'Zd6�l��]�<�Vl���r�T=�ՙ��4tF�[�0��=���6QKcR:ӻ��T}h��������nܪz�Z�ѝ��r*��Vɉ4 =�<�2t�E\�D�L��]H��DD�8�:�N�ԯg\�X��6��'�a��8�	�i�8��N�[U�����3��P�������̤Uuk���*TE
�L�>�)���(=�uE��T����� �P�tT05ޑCXlxVHYEB    a482     f408�t;d�s���tY��k��O�w:E�����>�
�~AM9�g�DjN��kJ}x�Y����ߧ�.�����o�B��g���`����Wb�_>�M��5�Ξ/��n��(��V��ʫ�V�(�`�ו��m��tw`͎�L�۹8P�I�-*0�a����04����FeU~�����=�@��_�Ed�������s��4�t��7�x.���^�G��<+��j�F�6ur���p.�\u���d��p����4H����1�8y��}���p��v�=�Ƶr�!�Ԣ�ѝ	o鳐����OY���~E�j�V!:�a�2���L{S.,�T&�'�TvW�˴���с���t�%f��+L�v~�]Z�>i� V�>�t�
b��L`�<����0�2 �d� � 5���JE�����+!n�e�eܭ=��`s�%>��QIF��7C����u(z�|�)��飳�?��T�L%�J��'��wG�}dq�����˩��{K�D���Uܞ֓��-��z��Y*Z��)���x��"�a�c�U(���qp2���,8��ղ:(�����ȱ�^�����mH�Ⱦvew1��<�%��C�eH_|5��	uޞ��n����]o�3����ų]Q�F4�c��_F�9�fo�vRU�(�
��y�J�}�X�*�����A�Ho��d����	��_���:;\c��"���]���穢'�}��m�	w�\��Ԇ��
��y�C�?����x'R����|�2$[-G�T��.]��@��3�������kr�$�����4�[�oe[EΓ��e˗�>D�[#Lz;�)
�"�e[�� %��Q�k�+o��+��c��NY�Ef9廮�6ߘs;�Q�& f����(>�O���y}̪�uhۥA1���GY�*�2Q'+Ty�1��jG�aj�V����ϩ��������i_��"���ت���i���8P��C"hMBHإ#�s�gp&@���=��~{��/j�����5]�����$S�~ZB!
ۈ�.=�2�\	ې�d���_�~�e�Wɷu5$|^=�c3�i	�K��c{��M��bY\L�϶`��$��k|�b���A�cva��4{I�_��F�ν��Q%L��.�~O���u@m��p^������1~^D�,�=�wT���m1L�4U���Lm��is��s�mH����z2t��'"w�} f��î���a�|C_����m��)�`�l��L͈���@�:�i��%��\��v��݀�0�-����(�s���K3�?�g�����ݻ�N�ŭ�E��Rs��+�[
nt�ebZ���uZm�����|�����ݘ#2*�#N}�ZH,1�
�לo�q��#vr	����̊�c�Il���j#�C��[��Xt�FJ��ܝ�w㎿:���tO�"4>-���K�'Z��Q~�.��߾�[Lۋ�BqA�f	�gC�6����[����MC�*�tLg�,��r��:�f!T�?A񊫗���ϻ�R[@��@\GQN�K"�M�^��%11L~���Cu�uS��\���
��� %��l(�=o�Iֈ�_0.�P�<O]��x������t�1��Q��2�erB8��o��=TYc̦*�^�#҅3n�2Z��1�'��n��/��[�q4�}2�P����@��{��k����~��C1U�S�鮝��:�`������q�� ����8�c��X�F
maJ	pp�̷��I9a=ʭ��qwgO/'�zN����<_�q�T�� ���o@�!��:��@������B;����˿-V���bA��h<�=���ߢ��s�)����P��_���;�n�Q-\Yoc@�jn�;B�r�B����{�%�bW�{�]r�Ԋ�Z���	Bc�%_k�?��S���+�٧��!rz��Mԇ�3�9M��E48��!�){z�\��#շ��b>,�j�v�b�t��+`];�9q�y�,ϊp�QɥNZB���;�3<��l5d;ſ�_���\<3�[�
b��.v�5݁@��/��L��S����Q�ID�W��L+a�����8��G�ʕ���㗶�܌��99\�����W&[��bj�[(���E����G�M����@�W�zK��ŎT<Ľ̿�N	���@564eb.;��$<(�J���3�O�Q��ò���?�)N���{�2l�D+FO�7
�u�x���m���5�c߸�̠�L0�ٱq���a|�jW��`B�� #u�G[�dD�Ō ��p�-���W��N����|p�ޜ�s�K�1F +'\��/x�G�O���!���ԉ�����&Q�ݯ})R	�M����1.{-�8���o�����Y��^��P�^č�W(�h�g��?��}"���Q����N���>N��-��R������7�@'���b�1��]2p-ď~�X�*`�$dp�*>����ұ��~w���%�I7X=4̍Y��i��5�V�.T~�D
w������Φ��f�XIH�ʒh��7s��J�]��R�y�"�b�>7N�w2��z.j�U)����g�(B\���`����d��.��y��~8U����F�3�<���/�"��0m�R��~����3o�Z�m��-�h��l`?�Z�M%�s۔Y��S���XK=��B.�_P��D�#������\�4/ў�G��^~�Q~�
�K�}A�;������Yr�@B���
���0�r��"L\�eۄ����@k=�8t�U��擓J��yv��8�]�kOB@���A	��x?������E����@&-]F�}`�z���`~	U�Ϟ;Y����&�S�� P��C�5Ӝ"��Ϧ�HUB�&� �ھ�F=�Ԛ��A�g}~
c�j�B�%�D��Ut{t�"N�������AVl�����o�d��� ��y�C�}����1&	G��ewE�L3������!5x0Ȑ �%�Sn+6%���	k[�c$��%�W�ɍcxʡD��V]S���n톜jL��Xw�`�U3�]׀�wuRá#�X���6�-n,{-����252�ы)*�>8�%D���+\��O��L���ߢB�lt?���5db�~�C�@'[�K��M��x[� ��M�����PTs�������0�P<��<��wi���x{��K��a�4p���23�p�����cnR&���p^aG�ꔵ+U\���������`	�2���G��|����v���wlm���[zKױ#�}�d\'#�p�M{�Ór��ӛ@����.��M��\W�S���rB��M��%�KJ<��@�����V�Q��y�0�������݈�_�% ��;�s@w�V�k�U��S�}��<^�1Y��P�}�6Xka�=I�[�zs����^9s��~+r��0������I���̈��7�ì�Es89~�����6��:�"��k��vj���m�Ae��bP3������L�3��t�����2O����{�X#���e+П��2�1kaL1�̗i��v1� �ԟx��V0w9�^<�&�h�i6ΰ�4D��IG:"b��CFtb�p�R�ѿa�ډ����rm,f��y!�w2���m�O�����}� K/���	�`=[�	='�uo��fܛ�&$禕PJ�	I�"�U��ٜ�W�}:m�
�V'�T�AX����	���\�Ld���Ȣ�M�pZ[]�������1��B��`�b�k"����ө{���۟K+e�����B]N�����`���;$�K�LBS�N��m