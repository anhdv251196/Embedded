XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��o�2���u?�o� �
ƚ[XX&5��q!��	�R�SM`�2�!*n$h��L����;��A��k�oj�;�|�v_��Ŧ�����#!1�=��:;�Ԑ��R�D�r@�Z׊��K���׍�� �������3����K�'n���If���թ*X��`����}��Z9D�p.���^�rA��2.i�L�MkL��+<�B�(�7�%&C��ڇ{ol��]�t�Q�)��A�(����B��{�l$�I�G�4 �i�o����*FTw�v�$/�Yt�!@�bw�÷R�t,��m�58X-�ȏ]7/��2���� ��țs������3�������&�3eF����߸��c��ZF����U�%Y�J���N
�>S�9S�I��ד��㤼��*�y��_��n��|�׽�S��֜�9��3҄u��!ݺhwu�CQ�O���1a���d"��6kd�ւ����߉̴�nW�V��������>H?T�6�;�@oP�,�s(4���X�p��SNգ��^��A{��]��3ۀ��eÞd�=�_����ߪ�%̀[c��e%�I�Vb%��<�=LQ�|�rk����ʉ�)��CB������YD7~� ��!$'�fO��zY,��4���6���v��K2���Й䠩���( �v��yn�K� �35�J�c�}ㄎ�x�����H��Q*�Den@�u����&L>ѕ��5�y�,U��~�#�XlxVHYEB    1d06     5c0�D��X��U�z�i��68[�~ �=7��x�՗]	wE�O�!d}0w�_|�?��Ug�جu�Y��|C@a�G��P���C}�>^�t�~�ˊv�h�6��}����� �����@����E���ԘX��R������`��-k�7ı}�	+b��g����}tǻ	DU��u"8�g@������Ѕ���a�4;lS�SWq�%�'�KEzXiA����j�;��F��+�m������A�ִ����|�g)�.�?�,�=��G�"�͟�ywi��3@(6��]ƥT.O�2HKE���5���A{�2�oCb��������9�^M�zt4�r��h[����RU�5��q&g��Go���
��g��G���� ݋`�9�˪,�|��4}���F�~>P��D-�[bD�i�*q��(�=Ծ�V�LC�����U���M�`����q���7��;�KMÜ7��1�����`[�`���U�/�qm[�ceO����iʡj3|
�1��<��(5�#��D1�&X�	$=�bz&o����5����v��`�<�{�S�H¶��pV��y+�lKا���}���c��mK_�+%OVx��+9�3��^�l[�5���ǖ�J:�jxF�8��O�U��F3�El)d����~�b�����MǍ؍�2��X�����H����E�!�C�h�+����_Α���	�aw�V�.�퓋~���bh��{�o�$~�1��d��D�/��Wت���*bR�.��e{�j�y�NI�ܢx����1�7��`���V���:t�,��R<]	DK������fv���E��e����L65e�g�;�FIA���1e��,)qD����/������d����mqa]м~d������ ���L6�H����/���I�RK-+���2���fzP{}�����G�w)��DT����BSȯ�,�-��'����E5�����<��~�t.�^�����ҤOH�Dn�O����-ȫ6`As�+��*�0z�p6w����:��<�Y���ȅ��ٙ ��z��AL< �f�k��j:�ɂP�ȬVA����b���D�g�j�V���m��,Z����SPul�p4�[�U��Y͙�٨"�Iz������O�/� k���ݺĠ���P�gj����2ߛ�������靫*4�^ ����F�iZ:³����w�n�1}Sb����A���mMX앂��C/��u�T_��Hr[F�7���"���,_��3�=�+�.Y�X�CC��J��ϫ���K�W��5�b�Ƃ���w��y��w���c�\�ԃ�߭�d������{2_DD_�T#�i���Y� 2kf`�oN괠��"�PZ�^��1a�������wp�� �����A��ؠ���P���*����Lw��ɭ&�bB*���G��