XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��LJ�3vĦ���d�������6izF���?.)l�5��j�X���a���x)���uK�����`P]9V��RQ��ז_y����nd�HΠ�t�ӌ���w�#Ү����M�n��q�2� �Rj�YV%c�T�-�l�	]���5Fӿ4M L@���i!M�uJZ�[�C��x���x�,�8}�T1,@8�fx���%�>��x�b�O-b�O�9-�T贵g�����z:���DX"x�~서9��b��C�k�Xmk�R�s����d��25�B�ݟ�c����/�)9(@p�M�]�kCq�l��T;~ͼ��W=ΒMIF������[: ��@}
ۙ����`���%rl	�YК�L�~��sw[�[�n"PFTfbzS�_�q��w�0�"��LQPE��^�䕲���:��_v �
T�F���/���tR�?WY��Hk+#�6!^j�����]�v��|���o�b!��X\`@����qo�
��پ<�q��U-��8�*U�#��/yPM��y�[<X��(^�n�����a%���O�?�ȴ��A��ft�m���<~�Q���F*_�M��7�����ӄ,`e��T�<���R��Pƿl��Y�:&PU��'4�9g���t�ڱOհ#��'�x�8#p�W�t͆(p�`��m���{����!���W�yz��t7M���\h��QT�+��>f]���݈��;]W7"X��.:�����ˁ�4��A *������Q���fXlxVHYEB    500d     be0G<��Y�5��g�<h�!��i$�zhZM/3q2�����%J�#'x�$k�Z
9
�v۵,�E�����ݸ(j��F��	���HJ��
���N+p��8�'ّ�_J�#�>���m#9�g�4��HW� @�<��?�;?��c᷉c:�g�V��H���{���%O��:�"qy~ Ui/l)β&��>u��#U?�}qa�[����Rh-�J��ǎ����7rB�y��9�f'�e�-�i�sٜ�������IjKF1zo=�y���m=�RxA�#1�b���xN�HI�gq��v5�v�nE�B}��N8tS�HK�����okȨQ2W_��JB~{-8�s�S�Xc�V#���deM �Z�M�FX�د��wP���{U܃�fbJ�.#��T��9��0P��N-��Lj�����y�z܍��_�ݡB
���hHP�T�A�*��W�YQ	�����kB���R�u.�:�ǌQ��̙�4-��7ah�ͣ�.7Ε�0����Y���� u� ��`�;���x艅�<���_B	��O���~�c!?w�2�q�3I�(w����:Z ��W�1H�a�º�.���
t.M��'�n)��;ca�iĪ���*����g�a�,*e���e��0i>�_��L`�~-u�Ae���A�Ģ�1���%���&�$?� �$�SB�� 
�نN��s�-�N��E>Y�@�y�'P�v�l�.�9���ݣ�ΘG���1�-ufC�D8�T�|]��߶�#G/-�˧���@���ڼm��4����.ˆ�!.8���)�,f9�ً���Zw�?K���ra]/y�j1�� ���ͅ=/�X��|ݫ���}k"j�GY(%i:�;¾d
����k=^��t���ަ�b�H^ILA��[�Ԉ�R���ƽ��.]��]֢ �������î*�>����h��ږ���2��۸(T�:)X�wST�{<��bN��?����'qC�� Mldhk����ʲ�=��P���{J��#�-i8�2����@��L��3G�>���&�݊���o��f�F�o2A���nW�w4�q��''Iƀ��t��w;0U��>X9�7�66����/a� ? [�I�w�Q��ց���_�m͐f<|A�Z[:���E\T	��U	{���U��P��poܔBb3.!����2��PsbR���5��cFB	뭪�=[����S������_��Yִ�?n��_[bG�?�=�,�դb�JI�uN8��q��'2�;�~..�����|�k�u�z�0�Ӹ��W_���Ru�ѕ�G�6�/_�����>;�`9����$OU>[��k#��X��N�����(��Gj�۰Mg��M��/������õ�>μH�\R
3���蔈h��紞���~*�AS�$�7HW��l�4�כ2��������^���8�9��	�r�o֦7"����C�z����/\,^�I	⭄ ��n
a��׊�F ZF&�k�<Ry�{*��, C^7�vE���Y��88qEZ���{�[Ą�)���Zi�f~'�%�*�ob�1}��R�`�4�+�J>���7��c#���GUmc}<|�2P{ۮ4�Ж��&U���h9�N4N�yT�!hI��J����ap�8�!]b���m� �_S�:���v������2*z�G���7x[6��#*�kx�6�ڲWق9h�̬���6Z���K�4y	�]=���R�������]��|�˂:��&s��%�X�H�@�<g�F��(��kP����FY\���=hvw�3�n�X�[�kw��3�����e�)�T� x�����a���Q��n��	,��
�)�D�cv�D�˳E��d����{H�4���٣���<,�4�5^�Q��Q�+^��Iz�8V3�t�"�/��O�aE�eX{f��M�F!�S{c?��IB뚐;��8�1�nr�|�@���H����%��pM��C��[�q��-�^�@����4&t���bh-14D��Reh��Dhx���(%V�t�[�1<uS8�M��ՠ�9�{s��Ex��0ON��`��$̙l�k���&%��d�j|�6����w	�@�cd��m�Е�Z�sAhr�pǳ��	�  +T8��Q(?}�i!P�i/0,U������>��-�Y��F`�(�w44f�yxi��ON���_�D�զ���#N��3A@n�A�&��[��O�>�X�)*�5�Yb��4��AY�UH{>�6�N��nI�WZ���� 7��X����fdD:Da�������R��V�V�ލ�[��%>5
h�d�t8�?Q�]��'����Ro�x������VLml��8Vk�D{�]��(����]
H�/����P���$$�FMMs<w�������y��B�?���<�����l�ۣ8��cn�!�6�7]w�0[+m"X�O�����_i�<�/R؊Օ1�v�f���ߺ�,��B-9,?-c�xo��ҧ̧.em�,�rd��p[��@4��t�O ����뻏i�[����N��>C&�bf�[�?	�2�+��
��
�,�*xe��OK9�M�ѣ���'t߈] 2�P
�G���{s�٧}nN:q^9�j+d���Kg�����V;��c�>��t�8�Cmu7'W���s����{x��G��o�����Z�� ����W�4Q 	WQ��.dq�����.F��N�
����K廖��+y鱑���A���SE)Y�5�
�W�0�Oe�pWG��T�l� �d�]�J�<����{�mʜ}Q�4��Y�e8��	 �7�"��x��g[y¾Xt����[��@]�$%�S����T=����p�.�?�7K�+@�O\������@|t�+HJf,RT�ה�׌D����"�3t��Fg �����=r=��Q�䟿o�|�f9S�_I�