XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��\��>@g?�MK���ϙ#�]�z�t�A��	?�<�/(lQa�PR�h��G`Bݶ��O�>�D�eE��j&͐~jpul��fg�Z�E
�������{z�"�O3�zm}�����oeM�/T��X9`gZ��QB�7{�K5 B��Kr̿�'U'�昗�
�4��b1H��wa�m���ϰV�A�8URԶ��9� �^��,�~�t�Hb
���=�l������'�$���bq�y�|g�x�홚8�x�h
]t�h8�$� .�guX�F�֕|J$Bj,�n�̃���x�@�bzx��=h�T�>����C��ɤ��l��B�q��jzmϿ�.:�p�3�D��+wGA�t"�@�.��G��O[��<��
��s�O�����ֱ�N(B�	q�)s!��E�2�h9b�bZ?d���YתT�_v�W'�Fv��-�Dc��z`aD~P�Ғ��gk"�	�*AVs�a>��M5Z����Ѕ22e���
�E�5���p)I4�C6ަ�c�#rh<_�eN�/���ؼ�%�8&Чƿ?�O�yo�v��������K"$^����D�x1oǠ��J��5��o$g�b$�`�cE�����{ȟ�GJ���!�ߕ-�x-�p��������������)]�"t�é�U���K(դ���-�sNw��4������2+0[�d�J�?ib�p��P�鸋��Ut]n}XmDhq}mU�q�f�E�@��xKv��B�MwT�XlxVHYEB    3a1b     d40�J�CB�5�6�4�Qr�������;�6s\�Q�n~�3fk��T:�z���*���Cە4K�Q���uA�Ky�h�3
F�m/0.0R�NX7g��^=���3�.]�Ye�Eki�ˋ(2_$�o(b9ף�7a��'4<�2����t�˾ 
�x����Cl��1�Z-*���I���-�X�?���ɧT�4mg������5'	���i����5hd�3H���WS,0B����@���4I�a�����PO/��dSLX��0�P ��*�aƂ�U@S�:Z������-���4�O����R�"�{��2\��u�ٽ2��*�.���s�ĩ��������~���;����:�w=�E	�*6�X�^�{��r�5�K܌��*��,((��Vh�E{�W��.oL'�5�o4�zRk��p�Iɞ�;R{WǃJ�w��N���Y;���/�������PS�=Ynuz�Ӄ?��N�p�wTs�V���)IC�Cl�	af�ηbѬ�Ҵ7��ϨkR��#�M��) 5�.}k�B.'f�W� i�f{K+��\����v��Zu�pD�#��Ñ3cZ� h��b6��O���?ˏ��o 3g
Ŧ|�?,k��S���*��7�'ڎ0��̨i��u=�3�k�E*���Aw0��D�%yk����9�_Z�љ>�\��c׼�A�4�wn����@��eK���u�'I��L2zP�8����b56jB�@�޷���U�EXYم6I\��K$Ii���&�U�"˦҄S�x?�Ki%�&ݫ��Y�ɭ���yJ����CP�gEH1�`���c�-$H��L)�������4j���^�yb��	�g;=9���*����*��h�s���Ȑ���Q�uq�S�=�K�ǯ%����[�l�쿱%���>�����,U���E�$B�r�QzW6���|�EU�l|*��(�y��X4�Jb��`����j8U�����k�K�t�^Ӯ���|��-Ҙ��kҝF?<����hS�O*�Xucs�1R@�w�����n��A�؀��,�Q~W:(�AB����`���A�U��n�`�5H�bx�r7_���f@;pN� ���_vD�^~/�˞���Qn �FI���#�yYc �����:��Y6FJU[*ĩ̈́4̄5�ѭ'���W��+]�|��;g�X&OI��I�󗌭|R$N��u�xx2/\V�����G\���_���4Il�F���ûC�+n<�&ɠ�v���됗�p�l��%�h��a��v�\��&�r��a,��z�Q]#��IRN��h%
tV{���+@v�_I�]Y�}7���#n'h���zgp��>
�E���5�_�o�_�j�F%K�ǒ�&2�C�R� �Z,�4�[��;��hq��1�Gb�?V�Ԕ0���,��Z�ĕ��XZ�HXaaTv����� ��!Ӛ��-�u�ɴW��
AX/ְ�.���Y�c6�JU��'��@j��e��Ɋ����q˲��hγ��>�-%UŲ��2�.A�{(��~;Uh����J������O���kn+I_�\/���RK�9m[jq�D&������v���mId����e#�U�и�&�#�*��Tgj�&�/GJ�{R�><V,���.D)�D��Ǧ���0�vF>g�,�,ygM�����z�����.��P���у�	�E<i���k���c[Y`�j́M��Y�ɕ�"�F���՟~�	x� H��V]�7�ɰ�y'c�e���ESG�e���k��$�kaL)D��|���QTâ��9�@|H��M��}����{j})�̍0��:�z�ey�c�б�Q0���R,L.ǭF'(���hLh=պ:��M{y.��D�se��s����{�M?��- �!HH��  sc�'��Ab"?;
�bV87k���^㊪b�Lѧ�ٻQ�!H�ݬ�p�7o�>�h�����F{ I�8�`�D��ڀ��o'p��p�¨%��>����		h��f>ޠ�4Q���4L3T�L 7�7d)���ʺ��$X�C�4)�l�V��r0߮�:��J-�c���s�!�Ww������2�^�Wה��J�{KG��ϗ���/�"O�y%�ֳ�Y�C�&q阧<N��*2Ww��Q�D*g�4^#u��`����>�(�>��V�=Oե�Ʀ�;:��S������hx�����1�j���	����pDy��b,5߶�ޑ\�o_g ��Gj�����Z{Y�Qm5�UWز=E�n�	�*�Y�8�.�;=�r��K�D@���{L�I�X)��F���Q����DLJw(��T<�:��ƗP���� ӆ����х����ͷKz]=al�~Hi���{6�w�]B�~,8/�l����@`�B���͹[��ȶK'Je9��צr�� �
X-��-�Ԇَ�����h���v�_W}�����j#��qg<cnN���z��4
.�}(�\	1�b�aȎcbI�3�ҴO���w6�[�X�~X1-fr^�d?���wyc�n�{��K�5.Jۛ��җ*����_�$�¥K�lx'����vH��8�9۠�i�7�M���&'�Mߥ�F�][+s��C��� ͤ�g� ��E��}ڣ
�I3Q���@���,����=2���� ���f�
)�ܞ��'�9�0�	��5��v�`��L��H�F�x՞���E���I��{L��CL���Z�a��c�s���fؚ���%����3�I��Z�8EPYV��@w��K2����m�A(3�ڞ+6��N�w<�b�h���y(�4&|p�Dy)OV�%%��O�M���-Ïb.�����G
µ�dAѠ-���g�0��}���>z��p?�k߬� v��n��/���	^�"��Kϴ�э�^����E':y�vJ��p2� ���ʩ�JKj��!]��P��W �j�&��E��i�4�ڥ��o�\;M���H�l��`����ā��!ڤQh%>����B���x~B����ȗ��n�iH&g:�x�K
W����5jj�Ҥ��taL����W�[�*�',�=�2.$)�l�|�:6%��<�7g���G=X���	�8	"�������8�5�S �s���K�jeƥ �6���eE�i��p1ueEW�J��(���r��,�&����n���TK�]D�x �$j�BF��d�?����٥��B��m�~C�{�NLn��6�Y�$9~x�)�	6� �~Dt�;��\�F��Li=�O��C��!���c��7l
�S���r