XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���F]B?��3���Hb@�aD���rS�^���g��I*��Δ��C.��<|Ä�͸���X��C��rr&U�t�1q����V�	6�z�L����>�ڙ,�_h��q�
�	R���4��3V�z���x��Y~:�VlGxY5M	 w�%G��pZj�K��O۟@<�f�C����Տ�ӻZ9p{M�K�0��-R�#dDB�uP�#L4���0, �����5X���9�Ā�'����A���l3���|C[ý߭x���9��$�R0�D~j2�sP�[[dĭw_c$u�D-�D��9ZZ����:<
wDr�IZ���h�|��,[��a�E���k�u9��� ��zw�g��94��C������
��
*î��.zEh� �=�%���ȯ� �Rj%~e?կ���?Пt�L�������f��l,�4�ݯ���AğKd=�(c/W��"ܾk�:�˲�-�b���i�h�$��a
��B}����s�:⠰�����s���%� �ɍ�)�$Ho5#�m6���%d��#��[���m~��k�{֏����Vp@Npkt�d�Ɏ�xĉ5�Wa%�d�]#���:�~(�����k�������^���9Dݗڴ��ĵ˂�3 ����q*�1te#ɟڿ�� d�q׀g��A�e�v�)KaW�eq��tB�'����J�������~����{�-zv�o�(�vj<}�����ы�%�2�/"��ŇƿyXlxVHYEB    3c92     900�KR�2��{_���hp��C~)eWE�͏�k��z�L���^ꑁ��Fl���
��~Q��;-G��I*7w�����PZ�;B냜���ߴ�k_�=�Cڕ�Du8��S��1����q*����M����P/y$�84!J�ʩ�c�Yd�ϓ���ӑ�dY�h>�r��}�}����|��q�7���0-y�/�d@ƪ��xC�HA�(���\�(��r~��v��mcT ���+��b�Tf��ۑ�I�W�L|�~��b9�(WG��.�o%�������>��!u�v�#2I��	K�v6J��={�y5��G�	 ��\ ��{AV��	x*�-�a�I��X� �x��L�+�"��%䰢��s�s��%V��%#��P�puo�#���Q��4���(�]��u��	��i�#B�����j����8��u���]���������	xg�y�"�-�a9-;�g������Qs]��W_��SS^��o��i'yK@�vΝ�ۃ�jhY���/���������a���n̨{�p{�����{��AY�&�"�M�vؐKS�KX��\Pz@B�$��
>��D?�F��l(Sˁ�ʠ �J�j�6&��hPt*t-E%�Vj+Ya������L�V�4f\�->-_I�/�ρi�8 �����Z��AJv���+�X�����y�P��5�pA<�j̸[�N=�U�(�ǃV!�6��r����S� �������cz{�#�lTc�"��]�pp�2�'�FH{8���&���
������?,tmd�c���P�/h�����u7:#�5�f钨%~�<���NB��N͓\�p�\A��ұD�w��j��z][��o4�R�b�RN�uk�}��P�UI��6	�wȕt(��R~��Z�%�f�TcK,?��g�����~�;%�;���ғl�F�� ^�L;jn��dw��k�"�[��������YV"m<��_&tu���������yS����K[�،�B�=��a�1V��Ȕ�����e�p��q�T����f�M�ʁ@�R�����'��x7�6�7t��1��Ƙ��xs=��!����~�l�>O���Բ����N�lLƓ`���?���T?x�?��&m/yg��)�E&=}�h�e)T�H�Դ����hn\�vB�B�^��m ��*Jݔ�/(��?g��j�^�9��_�8���>8U���G)Jzƾ�ԏAo^.��Õ���t������X�)��4�������Z'��W0,���K�龌$��xh�]�H����d�l}�����+d�U��5����&�TS�{�6�GΌ�GF��ߘU'&��|��)&±����#�_Ӽ%��g��j�w�Yrm~�+Kb� ��s��-V�G��P�fI�XR�煽rv4D��z��,��cN�������!b��q4._ڌ<#ۢ?iS�cp��XJIxU{�ߑ��Y4�8��+!�p<���U_�2ꦅ�)�o�.�C]t��aFI6��r��L��J,�������|k`�W�N����K�W��� B�{ `Aկ�I��t�.'���{��wt��cw�b�����G��!�1�
[6d=�.q^�Ae����6������b���+�~!G��Q��@G�ϡ�1�������`+\D���,�Ԭ����#a(��J��,����2}�}��%iQ6rK۠
ȓeqƊ(����H�Ќv���_�?����%��J*�[8И�eԢL�K��n?�Os�"}��j��.��F���/yoW�l2��%-3�(�:lJ�^2k-����u�KR�f�97 ͊b�	������rl߫E�ɛ~�j��)�J~�I�$Qw�5SM�d�(��T��R��]eS :H�jy���F�̫�؝��(zCS���=E��K&�J|:B�H<�S���|DH2�\�h�>%���H-�,��5������XE�DH�_(v���p���`������O����b�%1�a\RC̤g��wc<O��gݡ��}����I�1��z���u �,m`�k(O�\��߰�,�?�Vc
Vy4�ڴ����Q-�g��Vs=��ڌfF�>�o)�З}a�zK�1�� ��Ʌ�Q��-����<��;��ù	i(�sX|���<��#ҶMk���A:nЉV4�/o]-�e܀��Խ�*[�+ۤ|��\K\(�Ca�?��ſ'E�����uMg��l�8��n�n������R%����t��0�