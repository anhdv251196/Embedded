XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����{�=̹�q��&�G-K}0�#$��IE���um��/���g1�Fw*�����|C+{ۡ��?�j�3� ���y{��z��Ŗ���W��=�^�Z��L4_2�
�R���ք.G�E3/?i�!J��}!"k_$/(+e�Ɛ�?�qdm܋�ʩNe��S�CgaR�2��t��3�QW/����؝�L����}�Q� .��1�q���zY䧁��\���֛��?��J��]�R߼��-�Ri)�T1�F}����=f^��3� ��ُF��)�b��`J���Ē��JԔOGD �LV�O:8�����#_U(�=*�+Aeu����;à�}y~��-���
��I�-��@1r;�k��7a!�w'em��{�>����N��-/V��/�����)Yu�@	=1U���)�	;�J��b%F<)l��U���\��[��h��i�7:dQx� ��n��P��'y	OЈ���4�b�	%�/м��Ý��� �@�s�䱦�+�-�;��$? ��^ _�L�?ӲlႢh��������(Ѓ�k~�V�	Է�bsPy�v�_;�S��w�Z�g�}u��":��z�x��$���������Hdk?E��4c	����u��	2RO���6�frצXzVe����u/}���IX����������(���aUl��P��R<FSz���^���Ѥ�=�i����$_��#b�*1<���UM��=ڰ�ex�� �.aQ�K��`�XlxVHYEB    156b     590rI��B�7���y�m���i�Ll7���n�L<�JwI�L���"_k������G��Y�E�H�/T�=��|��s�Z�T�}<
����v�"~#C H����A�ej�=o\��V3]�g����	ڲ*��}F�V�,7�(�r>��x����%X8^Ȓ�8��O��ND��;em��hTO�f�8V`��_�mjK��#׽*X�����c�0����*8�L��7�a��N҇�@�D]́�?Ew�q�`C���1�ǥ�w��q�9�ӗ��ӭS�#�'�bW`ڶ5W���p]*õn�)X��=��,M��e���\���`�=�&��꿺U����t^�(����@O0e�ٲ~:l��^Dt��j=��X��<B�rm��s#��_yX�o�@����
�����{�@q���]De	�������~�&�>��2`�?�Ɏ�t'uôZ��2g~_0��{Q��ݚ����s��݃ԛ�Y�'L���Y(���BV��o�h��e�[���yM֖&�#��y�%҃�B�с_q��1Y����,z2���O��P։��;��_�De!��K����J��+�P��eg�tF��K�<
�?��_h��|��}my�9E�^>����l�#Q�ʘ,L��h�2)�p��k�y��Gd��]��ݼʒ�E�-�]Q=<�	�v��SɳN;����{�CW���!�$-�HE3�,�8���#'��#�*�_8��=I�C�I��[��a���ax�]����*)`�������iPJQ#f*���K����� an�W�d'D&��#p# ����.[���h� �l5���9��=�?6$����t#������%�ԃ1W�W��:(��9�Q�?������ri��A5�C�v^���Mf��.k�x�Ѿ꺙i��,y����ixC�vH�&���a�pp~׋����c�!����S�@������ː�"�X М���4wCZ�ٚ��u#����EA����H�8���u�Wǖh�+�EG�������-.���-4��X���b ;㰅;�ᛥ	'5#�g뱒f���}�t���7h��9����Ê�35�N����r����)�5��Si�w��\ƨjT����H����BZ�@�;���Fϔ<�6;��j� �P=�r�%6)"�Z	��n59�\���]���y���p����iq��,��{΁���CAD[�5��L��cۢ�ͽʦދa�ֹ`��� ��J��CG�a��U�+��@��#�"L�.pr
��-��*f�������W�G�������㥐z�P\��]A�J��P ���f8�0����_+J��ۇ�� ��h��zϊ���ܔ%x?ΕE�N�2����֝皪�
�IjR��5q#ZZ�s�R��