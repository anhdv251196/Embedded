XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��j��K:*L�Br�`
�h��B��u5�^+xCr�7�.(���5���C'��Fh%���]��	�����y�S��r��X�w�y�-E��n�+�L�{�����Z��D�Qw��/�<���2�� ��TLվ ��� u�W��h��"��5�S����}�C?�Օq#F<�_��ך5��3B�J���}n��pf�V�K�.\ϣ�+�}a#v�0� [�I}��F֐4���%��=b-a35?C8/���y �]<|�C�v��W,�6�ϕ��`��8�~�i�qB^���8����ȓ��B�ѸAHҦ�x��/aM�\<<���g7S�Ŀ�3&7�럇Y��}1�	"�Ҭr�(յ��H��'��"tP�^T��&0�p�����sm���kH|�6���p ���^��7�������y��I|%�a���C2��D/�Q�QB���zthn���ݪn%�ۧ�-˱�������_V`����M�T�$�;�O�OQ�DN�.���(m�ze�wB��%ì}uֿ6�!-�����<�<0{y�&��{���n)��{�*��2,\Қٚ�V(�f7�j TΆ�^ײ'��lFR3�3c뵄&���$z�{���}lN�*�8��uC���*c3��X����=9�*z��D��Z�zb���ӱ�m����O�j�S�\b�XoH���<�rǭ�Yuײ��*�u��c�͓��T-X�9�8HFsE�"�耶Q7.�۝�6EU.�iXlxVHYEB    6fc6     c30��
��_շQ��������U�;|��\��)�:��z��l���uL2��	+I�� @5�al�M�R.`�K��e�;!~ .��	�W�~��y�V
��si^2���͗Q�!h�Ï�Br��+oI����9ψa(��1��T�z�40{�}ihlL�M��S�P��ƿs�0dp����?��������[�W83��I՚�I����!��\��8�l3A-��"IO8z�&F�p���DR}�>K�"���t�2�d���^�0I�E����8�f5H8k�>C�6�鵣pD-T�&~�Q��.�j����z�P܂������Z�UC��e�)sǫhC�[�������F� �!Y�=Ϝ	��g��e@�u���;�	����P:�<�o��|�V*.Q3q�q�#�6�c�H�-��ؒ��z�ؙXvl��p�l�星�<L��9js�wQ)2N�&ͪ��am����ɍ��EY	���CB1�a��t|!��R�%X��BlE��(�n�~~Z���7��� CD��`w��9E;��=5�l��^��*��or�RW�	���v6��T9����齃
˽�[@��g�HP01ڇ%r��Ҋ]2�Zq���KJ).��^����]����pc�'^C��)�*�D2p��u�頚��n�QT*����7�+&���j!����v��"c)$}�������8�;�`�[P}�����!<�u�]��O�M�i^X��ޠ|*�b-2���-�����V�Ou���2����e�-���ۨu�����$́$�m�VǊ�ҬȢ40h�uO;uܬ�#M\^�fZ��e|9�R�Uʝ��}�{S/�ga��t��3��%�f|ce�?�̚[�:㶀tL�,��߁�M���ulO_����¼vT2G�j�ժQ�*zG�ؖ�y6&�=�O�S:�����'@�w^ι�8�X9k�+Q���d����"�6R߻y+�~D�7�������:jx�xG�M��f@�)�h�x�'r(7b���-p���a��*��������L1�4D��Z:*yz67E��g��+�h)Mf�3�Z��vn�^�gr*��H���ʀ�l�I2I7u��)�"),�=��$hw:��m3-P�6z�5b�S-�8�Y��N�1��F���~O��w*�{a��%���*����j:�E�@���[�5e����W	IL�[蜩��zͶ��Q�Љ$�|_w�w9� D^|���vM�fdg�[R+BM����k�a�D��I=�(I��c���7�}W%	I+Sy�_am�aМ�4��1���"Z����'�أg~cX�੆�9p	����~�}g�X�d��R ��C�������f��d��L�J�Ṣ��Q��}L�6��aD'�T�_w��˺��V$��W~��؏&?�7�r�o�b7?��%+�I	A�{q���r0�P�#�$FhT��xK��{K߆��J�b5��:�@�@)#a /����� $5��D�`�j:��M���M�'Q��h�di�&�l&ȷ� 9��$&�zYo~��"��Ѷ{0��_wv:�>�Q���R��y�H":��$s�� {q�)�AP�C}�R�CXSE�����]���B�������ʂ���&]���	�|ܔC��Ī��`�/ˆ�������ȧ+*b�+���-�Q��_���wt���q��fl��S�tLO�9���W� �0m��l�sK8,�=����t��+�F*�����#�c�P��C�`�Df�р8�ѱ��F�&g	Hm���� ����R�����|�V���Y�c�Ʃ�ltߑ�Y���1��$$b�[�d��n
�������e/V�F0�������`�l@1�C�hY0���p���L��s�-Ac�;t��s���+�����r�i�/SK|�d0P��܁#�(IbAT��D�;�/��[������d�
�v�z]�MR*�Θ�*�G�mL�z'�b���ц��1�]�@v>yXL�8�z���)��h��w����a��Fa'
t�o5�t�L��kg#�B}˓R�R�-������!F���J�D������T]�π�0�#�xe�lű>��r_�9�$z���#Z�KgI&g2�c�H�k>$ܞ�4�o��Ⱦ<�Zff�z��#��7���o�|�pkvG��=ن�-� K��������"�2 ���h�M@2�̜�\ܼ�@:ۙ�"���Y
˼�K��L����ذ��iGxT97g�nIa�{`�5TѲI�Q�d�mR�3R�3JI'6J����z�������2!~eV����u�/�ɁJ'��6�
�Z���$� A�2���ޡ�\B�[���x�- qp�}#� �����	��䵷>�Յm]�����4����-�2"uLcQ��譄X�qS��q6nɪF\���"�)e��6�W8J!^�]g�*שȂ/����������)��ýH�P�$JӍĲ�Ҡ"����R�攭� �/u�je�,�d���4d^�H��%_-�>2�9�F��W���������X�7�DQ2�����h�ۅ��	f�i{���|�g�q?�#��H������1���7L)e�݀4Q�-���ݺ �P���F��d�A�;Ej�0��_��v��UL�����QYI�`%L��1�ۋX���HuD;��g�:����jC�Ŕ�E�D��
|>X���5k���8��R�j�b3�xC�z5��$i��b���j�RD���7����D�I�0i�4QQ��v�>h��,�oBL\�/-gw���
����g8�Ƕ9��A���Ą����s�g�=?�=�<�?}��U~S1��V�_����	��r(^���wv�pY�*�o~֪0�Y�����2+a-0��G��:�:6�<H�n׮a�0w���'�}����1���@�I'&�y2w)���l�J���z�����u$�ǽeS�M�f��z �x�$�JBn����s����	Nm-����}w���*�캰K�2l;����J�x
��Qa�`�GZ���`��qdw����E�+M��D��-�p߈/7��"�G7��Q�S��K���