XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��0�*v���34�n8e{���=�E��$d�D�%h�燽Ttv��N K_<�4��T2��+C��!��K4sA���It�6�M��.�:��E�S��R����$�Y��3p[�7�?Zk����0�h.�]��"5�j2S���1�$��W:�Xb\,#�D���_����[�Ԯ̥��1_�f������2Ar�9�~Ik��D�KݶzW�f��kD�j ��'!8�,���y��˨2e��t����V���[����X��B� Nfa&���~PMg8����gZREL�v%�����"����d��׏�t�Cz#���no�v�U����&X�� ������S���S�#�I��p�v�h[�H_��,��R�:�TE9}�э�䬀ܹm_h��p��EI;e9?�Q�X� ���l���&<�@^bK�8��S��6�9B����8�C�۰vm+�ɍk#������3�q+e,=2�іZ�m�����Z����ڛ�dΊ�Z�)�N� -�ʺ���9�J�G�xOk��t�b��v��yv3m�|K����EnP����a�zϥ7N����L}i�+N�o��i���yX1��o"���x���b����.�����hA�a��dd�T�O��
��p�帊Q<�_���Ӯ�I�`�Ύ	��!���B�� �����4��_�	d��܈0�
�]�A�j/�୛�hf*�^�6�R�ͧ�	9p�|�6k�� p��=����A�VE����A��5I��9���eVVXlxVHYEB    4a98     e80�<8:�Fs�[��]�#��W���Ċ5������UL���&2�b�F��Q=#'�Q�TP�@�K��$�R���I��z����@�����Fx�J�vX�p8��T�k��!/-ki4���
�v}�讬wK�IJ��ԍ���6Q��r�ʿ�<wJX+����5�Af�IVht����d�/���x���Xa;GHR��%���p��^�=�y#���M�P�o���,�ͼJ�T����'k�*�3� K���ш[.�ݻ	ֈ�����~��|s�բ��o�1�+�\:�E;M~�7�!,ed	�ܟ��i#T�/�46�fOy�;��u��F&�dHId2o�9��S�;@0��eI�i�Q̧Qr�[�E�{Pw�;��Žރ|B#~���pv�@�]v��^������:���A�FH�7�'����M@晶G�j~H��:vRu�������c$���!	�c�H3��nF֫^g�.���{9ka�Y��oFwn�+�v̪8���	�<��Qܾk��S�*@�Ɂl�E�v6��x-����պ�Z�N�[��i�)<�c"?�4�d�Z
+�ޡ�޶��c�{����m/���磲���rrp�\�p�1�nΏ�@�}+�[�{���\%#�9��/���b��:��a�����Hb�����lM���o�!)�jc���f��]�����_�^j�x��]�a[���Z�	6qb	B�Q������:��d��r�/�d~����Ƽ�,��l"�㊐ة����X�KU������z�=KN�Ẁ,��0��/�o�g��X��_fxy�w�,�^)��������'��i+�c2^���E����k���7#��!^�ᖮ6�ʙ/� �$ W�Y5
�%�jÖ��9y)מ��v�9Rt�F��A ���.�`À�d��-�*Ǖ��-�e%��t�~:2���7�ڪ�?�U���JHQN��li�X~n����K���[&E�"G���Tq��;hMj��������e����,�a��B�B�~)*��X��(�Us���Gvj*�w|��j(M��DK	z��n����Hf#��0R��3f���8��AK�0�dy���z�I	�.@؜k�\��fyC�r��|��j�z�������/RZc_Ӫ&�v��}�T����R;�:��|@nrujZ"��(��0[��(8¸����!]�,���$��c�f�D*�I��^�8+����ל�}��z��)dt|�;�m3���ͳ�e��苇��zU��F�{�j��e{J����P�M�� (�Ԍiᐛ��kbH����
��q��#�W)+%�ă!�6UQ&���
�S7�Vы����B/ܧ��3Vd�҉��;�S߳�BVw���5�ݣdF�����H�}���ю6D��c,A;���c�U�%��o?���#~��1Nya���Y���e"�l|�L�g�'��*N�y\��b�^�)��_�rzz�Q�Y�m��D"X"�ι�$)���m�� �����;/[�U�T����˾g7����S�����
��<�oT�λE��16��@GPތuM窉�=M'ͣg�z��+���{�*r�$t�3�qU`�<�$��aq��ƌv��L��7�t��}F[��D[h<�O���!w ��Pl�:���Jl��X���\���x���յ����%�}�;����yy�Eu�Η��U&�t�I1�{Ύ�{D`����o��0�O�FS��i��#�;��sԳ|`�-��F�f��� m_*<����N���wj�1�8����3�~ϝ�?��ݓU'0�gj]����X��8ӣ�-�tMi2W��ؘRa:R��p�F��þ$�E���{wȱ*��T��#�����a�FMB&E�/�p����Je5�5�I���A#���m]��Npl�r�^2��!Y���̛ �Abb�/=����D�ƿ}u�1R�%��|����P2k�G�y�V(<K_GGL��w�8{��f��t�>Wa"�'f)�V���뭟�D�S��P�c���s3b���|�Q��xip�e�j�&��k����jQ��0�[��!��;�����1��_�qs��-�V�
`tx�3'�<&TMc��`E�A���IJ�w��RB3Z�[2i(�����K2W@�H8���2c��]�]u`?�b;��@��k���п�ܫRj���@\�q�n�ATE�2J�ȚG},2꼦ƝaAm�c/�,�R����Y�g���=T�s5��L��=�=�{��P�9������|�<��^��P���S��#>�	�5s�_�@?�%�|��=���Nr�����۷ 5m`���J~[�/=�hh�`�n����fP>��=w�,�kl\b����K�]&QΪՄ��_�Lef��2�9�{w���V5��d��D�oyk׊��`������]����{��F<~�Ӎ�l@���)#q�K�$�VT݅�mͯ�M����{��꠨��7�Ɯ��@+��8���ޔ��}R8=y��|~Rǉ���~�ðr�di6H2��� UgXn�'���4,5�H���>�J�:�(j�����$�n�.:�O��_?�6~O��ܻ$����x�ſ�m�����P%}�z��n�t]�(�@�Uu�����+���0������ʭ7S��6�O�^�pmh�!4���	x����kx�p�}yq�5��ua�`�c��8�^{`.��yKs�Ӄ���q2�'�|n �ͶS�nfL9;�;b��ѭ��h�4������Ҽ4�N+F�hW�h���z'��e"�;T��zS�Ue����Lj�r1��n|"^����n'��| ��]Fc�س�;˵��A~K�O��=dx-p�ʣJ�ʿԺ�%�4y�����,�VO܄F���o�&b��"�E�3�e��ʃ�ԑ;�~��Q"ďE�}xڎ׷�	�hs��wT{_����'��Z�	�x����Ԭ\�fL)I�:bc-+��nРޭ�ud����*C=3���m����L/�����* T��@�=a��(� �����|7�L�$pBT���E�\�H��	�Wk]�������LR�G�t]=��6�����HP�qe4�ۏ�O>�ĺrÖ�<?^�	g�[da(�l띑`��q��
$|��a4����.2:^��e�J�!�VO>��Ǥ�]�ŭo��T�fÑ���h-��R�@��4�8���:� �U�{J=�N��{fV�Ú�����b���r�;[ϰ������T�-�2��,`/T��'8X�t.ᝆ��3�U���?!m���P��eĎ�7 �m�;�Ҏ��ݷ[� ���os��;���5,� (�8�}>��zfh2�K�kz'�$^�Ap[��@�l���B��"^C�w1�I�UA�-�J������I��p:�S�[�x��ͻ�w���LD���1�\���c\k@���o�΢pO�Xb��'�Œ��ye<g�Z_�y�bQ|�b��L�r���"I��
�טӢ8]=��ڢƹ��P���k����j!CD����&�QVJ�P\	E7�(F?�܌˦�̜!��}_�{7�n�/wd��̦ ��pg�5Г�4��v�9����~Q),�OZfͭ���)�(���,�@�,n|�cQ,��	!n�l�����r/�t��=