XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��	k
6��bK	��� r��ۗ�e��ƙ�B��U�mp��In;����١Or}&��ښ'�̛c)'!σ/�K��$.oB�a��ק�c��ChT~��ξ2�8D���>z��j��T����38e���dЍ��i�}��#�KU��n�%�E�]g�LYR^Z��>�8��i�'a�iz���Kvz��F"�tF ������@X����ԏ9f?&
�lK�h:8P ��ʇ�0�(�'�,��ܘ~h���&�<e#iI��4Ց�(&`zm�5-	��J~��Y��/&G@
�a�x��d,� @��\�ߎ��~�7{e7�p�pZ�Ne����P��%�&�!�a?��yӜUR�����5��:!�jZ��$ф�V+���Uhm���|6e.�����e��I�������i�b�Uj�}����IT���T�̺�N5�z�k�Ra�Rn��r��e{��X��'�Ҡ�i�Ԉg�ik��ɍ�Ĭ��� �i��DX����뵞:g��eG<v0濶���`��l{�Y.���U������΄$�O�i��@��%�_�έu���QDM�)��9���|m�(Ew?q��u ��ٛ$н���M7!�t���vo��u�M܃���t�<�뗊I��=�0S�tA�?,!a��� ����?|�;��n~��$З�s�}��g�
��bx��O����$� �|����3��*=,I�d��������K��JFI�#�"�T�й��"XlxVHYEB    225f     610���.���U6�u�_3�ύ7�@�.Rx_�:I��53�@�P�v0u1=~��a�)[��=E U�_E�TK$�flB
�a�6��|�3(`���dU�u��,Q>Ǖ�}J>���!j��h�D���f��犻]�'R��!2ZV�\�V����E����f�Z�!:�Q'�~-s��hrl�I������̨	B��I̎��+�f-��}�n%+�7eH��O��IՉ�Զ�j,.�r]�^*�0�i�1�Յ�RL�5Ȧ�Lw$&�:�����X,��Ų��3��6zjr�\��>�"�,��������-��jLhҺ��$�2]c�e5�f��סqJ~6��ݮ��#iB+��`u5�h=z��;���[^5�p�0�}����d���2.��e�T6�2�����liu��+ʝ}s�
y	O�>Z�yj.i�LںU�*�+�Y�� ���uK�	�!$��A`�����%�V#.�Q����u����}���2y���K׾��B�q\���#�J�%��m�4�Ĩ�6Ż�_�t8b�����"�l���]��9�@�qK[�B���~����8�Q.u�חٔ~��[��X>�F7�L|�x��\��|��`*:��po�=µ�,�#��\�]hq}�x��0է`$�JTy2��Z苡�R���^�����(	Y(�p����j�X��#�nm:�2*G������RBq��n'*x㎦$޽�P�������:c����fÉ��	Ir�ܢc�rHI�]̥M�Wp&�ܘm&6�!*`�hG�^5�j7^Q%�>�7�iR�=��
��}D���� _$N����DT�7d�+��C�@-œu�5���I�� ��A��~��$�`4�S�!I�!�g��q��]�/�Ա
��7[�yayr�6'd(�ѹ�őo�1=�9JG��x��rŅ�_�)�AT��Y���;W��c%�sJP��IiV߿��kA�������z�L�Om~f|u��ʲ��ҟ���u㏷R��������b��>ʔ#r��T��ץ�w#��7a���aK�炕"y,��)ˡ�M�WH�z�G����HN<q�i.��:&B�z!�"U�9��	�:�h%Arǯ����I�;,���O�pp�0mM҉��Y��/mE�եO6�i�)7�y���q�|�O�/��<��%���Y��	'١[Y"N�Y��,#}!_yY�⬛L[�V�
Л��-Sd��H��.uE����c�1P�.P]�E
�W⨲a!��g��`�zu���]��m��
�:�f�3ҲT�\(���%>���{V��^FKp��&�o�X��Bl�Y�	�_a�fⶢ�g:�����6�j������v�M�7�ֈ��#F�N�TP8��8҈�r�/����]��v�+���,>�B�y���RL�P�;�@��5t�ް����Ee�@.����zh����e�Ah�ز�)�h��x�i���]�f�ͣ�[}�1�)���Ш&{X���DP]�/a��}8"�H�^�/��