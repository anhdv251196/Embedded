XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��D�Z�<�2բ�}�W�1^,���������D�I���䣃Y���ƻ��0l~n�+'�?��ؒ��w�.9�n�� `u0�����glh�ݨ�I�Md�-�Z���C�Y���j.������śK�
j GI�lA�a�#_��s�42I ���(.H幒��6�-m4XG�h�3� ���K����M,��lO[����� e���k��D:�E渘�^��8�j�c[�<�#h�_�p�L�8i�3�(�j�� ���T~�}d�a.�z�%��ƥM?�ZrbBv�����ýS�Hp��xp"�o���>��P.X#�:�!Ȉ����3���~���HCy�l��C���5�JL��Ѩ�yg�<�	�b��0זt��uO-,���x�f�w��;��A� ��L=X4����姃��q�Z��܃Df���v�M�z�Гe\0Ũ!X���R�lb�'�i ��.pP~%е�nUպ{�]`)}1oAS_��vykf;��~�)biOSe'��L�P_0��]�	��L'��Q�h��3B~Yk-A�@�����PM�v�=�C(�����)�ZًI��p�|��SJO1f��t�Jҝ�z�,���c�ĩj"�쓶>6�耖���:#��&��/x�6�NF��j����P��%�����f/B��IyRхU���~
)%��0�
�Pm����[�?_2��x Ll���;��������}�\�&��X��1���k_�����ȓ<Fc��'t�����㽸�MqhWXlxVHYEB     99f     360��:�Q�[����D5��1�\wH��X���}�Lt'b�jq~K\��p<r���V'N�]xt$�;\L��	�<�OI���Z�� �Yv�Cj\4�C��e�}]K :�i��8�Nmt�eQA�1��.��[���nznN�i�=��^�)�W*"�:g�9
t��%mL�\�&�/7��Y���ނq����q9��D \\���w
�ua�F�#/*h;:7!/@��J^-�/�E��e�F�>
j�����YJy>����5�e��]��d���M/g�@dm�M��~�Dd�^�4��5��� �A���ꁋ'e"s������L	��~k���|b��,�[��t��1��o�6-K���L�����������Ӳ�Wy��3{f�3F�fǜt��Sz��=�C�@A��f�)��0س4��bR0lf�L�i0O�W�e�����K< �n`^�q
��Aގ��b�ҟ���|���}��U��p��T��^m>�
��N�cl@�a���T{���d5μk���
�( 1�c�1%��D�B�(-@�[?� Hx��A�����h�����{�Y����0T�+�:Xt� ��~��[���y>���fI'3H ��+2<-O��I��պ��?��抲���.����7��)��.|'��)�&��JX�w�S�����k�_�4�Ma'�=����C2�-���Z��� ��K7��9���K����q�.�d��3�?�zF�v���KA��\�vy�z��e���#��OE�I������i�LM��5"P^�C���׺6���k&���Hm��cC�Q��a1�D�'&2��^d����