XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ocF��+��&_)��~Y�f$P�p{���\j��_u�c+eu�Q��f����%�Iw�ZaM1�YEj_�;IG�;�.w����d����ի4�e\D۴����G35�*��".!@��!�R�gƙb�vn�]36�Z-�ԡ#��Ebw�x��g'7v�"ξ�	�[�L����� ��0	E(4��>�3
o�.QRQ|�;�x0�u��/�,9���}�v����&b.��� +�J���L}�%F�D�1�t�w����Kv���P�9�3�X$�� ��0Żԧ����Ǻ� O���؛�mQ�;0b��Ѭ'E��� 6R\��׷��Τ�J����c���1��I{�o-��uQ&=���q|�L���L_X�;�����jHn涀[Iݢ�,��$�~|$����@�fGG����@27.��c��2dQ؜�TB��c�m=�KB�n'� A�%�FcQc��M�9��֯���bk����XU���sK���������)��������ܶI�2-td�Z?Z���zu�����:�x��zU����	��?���Bx��qj��
�P�V{��		��k�3�r���4�p��ݢ���q��
���g��C��B!�<�?��$e�n�ɏ�EۆS���1����<j�4�X���UzzP74�W���m>�S������[�����$�'�����(N}�w�yQ�����H`Y�А�b�*�
�0i
T�54�S���w��y��G2�
��XlxVHYEB    41cf     c40�yMSFp�۲L�����f�H��E��\٨}���{��{v�:��d���bRUr�/�����Z
rw�K�T�jO���י���H��5��r#^�{#gYo�lzhU�P��⾚ˮ[7ԭ�I�'�j�O�#O#@盉�*�}�9�܄C�X��D�M�KbƁ��D������% JP����̿s�!��&eZ^'p�o�<��;mB�Yd�汻~ĩ'X����Z�&j����ˏ��Vs�r���+=H���7&"�'�]�Y��ZYl�W���>���GD�{]"�h�FѺW�Uh5Ԗ�G%��)$R�f�R�v��ڴ,�]�Co���>3.��..��C�"1�:�t�5���[ۛ2w�?��$>�َyu���-Pf��HV�o:�
a��>���-��{����k��Yz>`1��]�/!��lEltv�г�O��>x>gOZ+q��G �Mm����^[)V�n*�V���F�X��i��8�MAV�����B40Y���>�� ����g���^,�k9��(n�����uĻ���(dݵ�S��+�����X��U�0� .Q����ܼ.� z�)����?�gP0_UB������{f�V��^!o�PqU�A�0��b�{�8�2\T���?Zm��}2X�.��tO��E�²f��j�d��y�D8vBN�Bn�N��㣝Ks���O*��v8̕�`���kg�3\��K�*��`乃9�
��2�b<%�`��j���:���2rAJ�G��3E(�r�U��&�~>����<��$�>z����0W_�D[�-칂��7	˷�`V[:�d`�^��@=W2<�����!6$�������X;[����F�cUTѢ:U�E���<��7*嫁��CZf�S W6�H##�b��۩�����΋�/�WT���,�W+ԡڼ\p��U��TG��F���Sɜ��
�{��|az'�X4F��AeB��e�ܥ��ϕ2�Ƹi�,/<OLD�qs��~����5�tF:�ߕ�B����wE3aG0D�N@

��Z,'�f.��#�A���(k(!oS7_�%v��ٻ��@��6�_�0���x�o�gy&x�R�Xg&pSu�v�Lh29���ϳM�B���"j㤙��T�1��*��`C�&��窓�+A���C艼����I�?��<FT�J_�~ ���H`�Xp������R+sE��:��iO���v��\D�C�7h�zQ�9�D����^��v����+XZ�ő�x�߾��ټ\�����!���� C����>/�����-U��Q&�a�Ci��K��l�y	��B�h���Լ��u�)�ί����(��m�jXv+���,3�}{Ϲj��'�W�a��h�裁7ŕF��^�bM��2�h��' ��%����R"+wY��;��KǎJ�cRՊ�oc�{DHI���IPc(M/za��%�{���[�t��J�wi�%�Л}k�$�Vmr��������|2g���{���n"�F�����UN�n��������j:O-	`O�U���t�r�,�[�E2���U�
��멖a��؃ﳖ�8`w��%����1_�nH���	b���RG���p)�)%Xu��,��F��T}���y��M�1��H�c`��4�@�Ed7^��,���6\d�O��&G�j�+���e�Y�V�S�P�
6�.ܑ�nt�ˊ���_��(�� �}l�uqK<ӌ����k�A)d�T���� �ƫzV~��+PǚJ�����dS"5F�5VL%�<óys��.�����!��3!��N���H�Y����dʊWX�������x�Ľ87jAФː1�_]fc���`1�wF�t����&��8-`�5����VT	����egl<,~���n��C��Y��[��>Õ�+<�B�z�Ɉ-�}��J�� O����� �T	q�'��u��P��3�	[2�Un�)�����	�m�+b�Ǎja�K�ɑy�<���_ȿ� ��'8�������ߨ�G�4\�vbHvM��7Sg�y(Z�A%�I�w��񐬌���і�����P�g�Jcd�jX�erH}(��L�/Kf�gn8��ڵ��ܼ�ɗ!tϴȠ���GpVPQ4�M�EȗNI�\���({�$�i]N��-��2_`u�QO��H�?yQ[��ߦ�G�g�[��蠜�j��&�(îEi���a-г9lo9u�(u�&�U�I���H!RP�K7���]-eW+s>���w���p���N>�q��bR�y؂y�K�q��x
�@�����a�g�TD��)�t���%���]��Gj�Nzh���ϔҨZ�h��1�E�l�_y~r�tU$�����t�G~���E�JwrR0��4�<f]��(�W1�/�J�`���M�f����I%�I�����Ґt�z��r޲�d`/Yf�����R�S�ǈ�ԞA<��T�&�.�ʸ�b!R-���2�\�7�h���W�H�EL����W���O-9��u���a��uU I�nvkr��B�Y �
˪B�#{ ���)j2�'M"��7����&W��DS'�b����K�6��c���� �Z�f�6�����{K�!�ՌК]��B��1·��$!������w���{o KʺYZD``�ϲ��)�	��4��mO$!H�p?�)��d �?��Jd�Īx���gvH��|L��ISˣ.�{o�ʀ����]�s9����(%��a7iƺ�ph?�����-t��\�m�M�N�q�v;�	��#l���֞��YEƃ�pn������`��;���4XY4q���}��}�F|���s�Ba )m�_F#�:�m
!��"�<@��
���2��FcF�1�ߧHgy��3(:���ؙv���hG��q��V�/A�26Z���%m/~<���*����� Li�$x�*��Z杴��H��ӟrC��<i�|�\E��Wb�Ub�B�k����N��>�j�|p<T#w�E3ou4����|��	����ʠ��[�:V�0�.:0�ܔ{f_!ƻ��i��~6<N�FM��%ޫxS����g:��]��x�������Ǽ�B