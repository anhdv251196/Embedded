XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��D�9�.eZ�N��X�T'%`~�`(Zs���뺢f�jO9����IN5d�$�_��"o��*��癥X16]�6�����yΝ%����2{	� S�������������y�0s�$�k������ZݸG'��K?鹌�Cߎt���Lwȩ�+N�`oq�:��[�r(=RC��S�*�hN�?��_g�+$��`��<�i���_����������mh���̎���C_@����^��	�����\�ڄ?�ܴ �P��8�n�Yи�} �0�ɇuNvi�����>w�&[��0]�o����W1Lo�%����ϓ���?p�C@�������~��6o�*�ָN6 ۽�@&�n��I�4^��AS�Ox`��cm���U�M��F��4z����'6o槇{͌�gxE����n�:�SۘdӦ{/(	I��Sڧ#�����m!7�PN~I��葷h����ǀ/���U�^]��ԒuqY��o�s�b�1@؆a�͉E�7�d<��7¼%�YX�p�9�#̔@$��ud?
cӴ��Wr ��t+�;�hL6m��f)�YVe�/y�u~9Ѹ�(e^X7\���Cj��:���BvODR��%�g#�\�;�>�	ݝ۫�7V��ePɃ�Wo5�Z4�f瑧	.�9b�Z̃��yZ+xp=𵐴�k�ԋ�Ie�;���Y��ɰ}�K\���7�#�Z-���蒛JS҉.:�@*���f�7`�`�*���P��Aq^�*�/����r�!�Km�*й�&XlxVHYEB    1044     4a0\`vsst�}\�n�|��i ���ɖ���&X�=�
~2���v�'N�ۣ�+pP6��3�*=|v���}4� O�{ݮ�H�r�՛�j=S�(P���ZۼV��:�Z^���8�7�jMFLMh�J�uс/3/_�U7q�d`㢈uU\V�b�j4�P�E��w����~t����p�6�4���QV��l*��{|(���9�f�jx����'���C���!(F����9�.�p��<=֑���Wy6�%]}��,�k�Jڋ�����}���눧_�+��T$�`���F����Dq0"�� �@tR�66Ŭޏ��K8;��0�Ȁ�7�|�G�M�~[M#Hov��#��R�ؚ�݃����,Qj���̦]�{N(Seē���
N�؃B�訧�	�}M�T��.�`\A=\��3AQ�����Y����p]�I�Hk���ږ?6ŦN^�dj,��/ÝS0�e%���%��o����.�˙��L��@7\����p.[�Zs�kTœ����ɑ%?�b��t���@J�嫜��vV���6kT�!1c��j������W��h�=a;�ۘtq���q��J/%�A��Y��W굩`��1�����u�2Mg�L,�&u,#���8C��UԊ9&'Q˳v�E/O���KT���.t�֡�qw�:�uh������<gN��>���Ob ?��5'8�2Zlmr��J���	3OX�SD�V��\��j���t	ɼyTo7QX20ij2W���%s�g�ꑡ6,y^�Y�P@*]	yrD��px����j��8X���c���"����c����n%����e�D>�4��?�ć�< �=>�.�o�R�Є���UC��a<ǚb5.] 
k��T��[�fT%��C��T���i�0�Ц̺�����%ҸSm�g<j�W%4I=깢�6t�Fi/#� ���K�,׺����W���z{�0�A���R��k�F�R\�vE ���Sg���J��\�X�~.4m}Ag�Yp�JC�r9	����f��~�Tf�	b�2H��!Ò���zYa��CB%6?�A'�+���C|�R����p�#$K�0i�^~D�s�����y�s�-���_��GA�?1=J�+��a��4���=�)�#