XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��B��I��b���|����{^hM���~�ME�z�"����Q��Υ���a&n�^�#���:���nZ�c�������
�3�AnAԅ�L�TB���dE��w].�27�W$8�x�Ҽo�)t�eDC��~w.�),)�@]�E���u��RG��43������Л�Ì6�Aa���~�������~i�a�<��n5���/T�%�" �FѴ-�aS���I�h�;����V*C�ü�.m���;8 e'$�-x�H8f�������>!���D	�e����ՆȀF�]t~
E�>�9�%tQ�r������L>��#q>�n�[>�׭���~	��d#�����u�Rδ�a���Lg��H�ma����q�z��B�hA�R"vÀ��4�L3�X���V{1-���'�Y�t�m��-/=/��?5l���nV������o��b��Z��� �N�z����ʈ��M<��9Hb�W
̝a�}F� I0㢍͹L���4�f�k%X���h�@~�����,V�iJ���)������Cs�d��1[�q5�׬��$��7v~i$�������q���ؿ��ʐ���PC�hA�W!9�)!�\B.U'��p$Tq��5�5�r܎A�qeQx�.w|_!��ڌ�n_E���Bd�ȃ���tJ��4��|�t"Ђ��{`/��v��Zȝ��3���u_.�$f���lPg}m���<"�=	c}��񠛞�OMWԲ:D�2��{�6Q�3֗���{��u1�O.�XlxVHYEB    152e     580��tJƻ��׵�2^�U�e�mD�����K��&ӄl�@��Τ|�l����X�������N^�L��ƅ���t��P�������mF����ͥ� ��U��K^��rzL�^���N�U������:(�p��_�n�M��ݰ�~(����Ud�!���y@�LQw�hL0 X�Vh���v�VQ���/rZ�9~�ыT��1>�%*��;�N�M�d��	]�#�(���~�e�{wJ�l�>(��_��F����xݷ����>�o�s�ӅfCT�ǝ���oy� �� �YeÜ�[*#�=Eo������>�m2�$�$',ky�,3�܈�`Y%���4�*��y@����#�q��IT�
F5�hJ;�=�a2���2ĸ|���G�k'F����Y��t�.��P�*�V:��8|-
`ۡ�:��Lw�z��Y�h�݆@GŰ�J�R3�����XCx��S�盍��>�{�J�H�	��{c��e��TE��Od|���%1k 	]�6��7���0N��D��j������Ͱԛυ��kk[��v�؀��	A%d�P�o�u������P��L�
�+k���/�H5�`�s�:�y��ʢ�X��(�/Ew�	��ag"�5*`���o�|���0+�xB�V��i��^�|jlkòm��G���~����ꔫ������}o���������T�M6�����挄�C���l)�.���]H(�*����=E���2M�=�>pN� _o�����ϥ7��� p��Sy�i<��5���M\�IKэ6�L{ޝ��
������Ų��^rH�ح��18J�I��өM]��5�H���t�R��I�v��:�Rt�*Vq��^��Lr�gE������_���(5������{��-q뿭?��cB
��⻣�IUY�̮���o�P��]_�J2� %z���t�鱎�-,�A�h�u�ķ�#L��.PH���\Oe!����+'}E]/�W�D�*uV_�;_���!�Jv+���眞�u�<B�LgP�n�M��t��W�w�Tc_-<���iy���fI�.G�tHC��Y�7J�b���g{vO�]�7��Ke���1zkb�l���|)���L�KWZ��l��/R�L�!C�"�2�0&�*�I���2V��}'�>��9w�x���]��Ji|���K_�%;�� <�	�*9�K����]�$�KGk^��9L%} ���t���4�~��ޤ�y�sqЮ��gGF͉�a��L��זv��I8�Jv��6S9F�x��j��rYDz�O9��t�����ˏrW{�.�Fu	"�Q�D�`�p�&�D@A����2
�(�#͛'A3u{��!��0'��X;��