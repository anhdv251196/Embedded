XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����p}��P�AA���Wm�ȁ�ƅ���?!_2��J�p"����Ĕ;̫v���D��:'��g5�5��:;@ �z��("Qڐ'��|�(c�Y��I���q��R������/�9~-��p���=n�K����ɸu��Qn4Ȩ�s{�\�}����ޱa�z�xS� c��NI�x��a�������?i�]j��9��t�_8;wݿs��?�}C��ػmDE��W�7js�VP�l�Hro�טE�K���cZ�������+�P��QMt]&}��S	���g��cwxo$�n���@ý)�k�- ��t�%�U�O� 3"'{�Z}o�ޝv��4� ��6&Y�CƵ3� [u�p!�ȴ�Zs�Lꭀ�ʧ�#;��PEaIo9�����jЯ�q�%s��z���@-t��N�R���)��)X��H�5�[Ab��(�����F�&$�L�[�
?;�)�e��脾�z>�P�[X{a�R�a�ЋUS0���4~
nX(����C7�jN6Nc�'�`�՝�=]J����}�Si��`l)��:�Eh����P�j8�;M��wsj�͓OS����Х2�,���Y��-p"�>�[�߯Ld#+1^HB��pJ�A/��)��>e+� �Ғp��F�1:\�T���m�?Xͮ���1Q��yH�b5�+�Jbg������I��^$���
�L#�{zh6�<��~�<WY/���ҋ����eݾ��������~ނup���XlxVHYEB    156c     590���4 n�2��:�e5��,�`��R���r6�L�s�s\&Eq֪U��A�����olrn:oå9��4s���^�u$�`�.fѵP��J�'i˴H�NT�:�I4Hu�m�q���q5��wy�y�kG�F��l�8���(Yh�J��o�z2OD�\�,SJC֑p�;����I�f��S��T�#����Ў�.)�'zW���OvԶ�:T�����|G���*Ӎ~gS�i!�G��X�g��]���Q|F��W/����ܵ>��~�D@���2/��YZ��_$R�k{���E4��-���:��J�q -M�k��8����hMn����P�x���T,���sЭ?��Ƕ�UY	�·wU�J*=��/�/��ɐ~=���Uٍ�"�)�\ܹKa���`A8���i��'x�`�t��`�۳���G�}[q�o�k�A����	<��YK�n�<�h)/u"����	EU',5<s�����ѽ�rIt���}����Z�bi�)n����Ƣ���\>���cͱ��;�@���/k��'���m�0�U-f/2m����|	�4�B�edM 7�_\e��7�!�G���Z��X��}4�ls<|V�������ß����af����:itv���x�ӄ��d<�Q���g��	�0k��=(Gb�	%8�I ���;~��(岴{N}h�ʐ�=����ogFW53������=�I�,��El��k����fAyt�yJ�>Gl���D{�0�Vy�D���XՌU��ƺ� �9��<-E�4���?�ع�F������@�B��}%�	�����T�'�}U�='��k~�E�����)�;�H�����Ơn��`G��?CT��k������ʼ�/>��,q3z{�P�I��>�9:HF�[K>瀤{��#q���<S�g8�h��V���׋`���WY$�|Q��=nx��X}Dׄ}�G�[�گ+4Y���M�������yq�o��p���CzJ,5D�)�s���|�-h�2/6��t>���Z���Y���a h��c�e0*�W3]"�v�$AK�ߢӑ䋌�R���v��AD�V��-RMx~�8�4=�RA&����$���	T��|+��r0�>��# ��{BG�l�D�����bf˃^��s�qe����a���T2��aPG�\i��������6M ��29�^�79QPq�	�B�6��X�&�wg)��zů��<Y��/�}/]{�h��P���K�ŜVSr�Yi����	'fZ�@���t�� �=�w蠰ɟ?��l�t�/r��+�D������M�䎂�H�����P1ʢ
�d����~zJ�Wެ�q������3�u��١������AG{��������