XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ޕ��6��4d�E\�j�@�^�e��m��[��-�	HR�����8ǋЙ2ͳ3��G�`��,Ջ��"E��\`E�PE��ݹ�s%��{�b��Z�܄p9\�مq�}W��+:,�E�u/��9=il�q�p>�U�	���dX�iU���� �$�����(b��%���!�y��r�yQ	�n�@5u�i��J�C����Њdo�K�$�5l���ϰ�0���� �\c���[��ᓮ��a<��	)/��#k��0-��{���<���j	b6N��Ho���Px���VE�|�Q� ���8��l��Mi���«_/T?��D�)�Ŵ�	��wA�_o�+�j��rX����do�c������-	��(�v>P�.Հ��Z��/,�����ʨ�'+�-�Psj�s*��t�\�N�`�"��U�(��j
0�٥.�Z��T���|4\g�	���i:�W�)�rU� )���F��}x]h��'~�2F��J�{�!�����)��	�Rk���DLz-��$v<M&e�/Jl��u�����:�'%s��d�g�iB� #�Mۛ�ܞ	f^g�ZaL�;�#�Ѹ|FJ��_kF�2IpT���D�J����x6D�w�X�N0�D��P������j�ݯ�I�Ή�7�y�f��	����ܵ�IL�`��\�I�r��[���9a�l�s�X+�ȿ�ͻ�� 9�K}QW�(v�x6���a��:ř�8�����m~�{�6X����7����AXlxVHYEB    cc3b    16b0��ۻ�yc|p��Q,�/Ǚ=����@�~,>���*�����3��Xr�.����<��� l=Ǟ)���xu��� �p�My
��v�H�W$ǆ�`�P�}�x鰘:��x���U�f^N?`(��0�y������-��h��πU*�~̈b��z�F����7b�'��v���X=��>�}eD�{��Է�w������ɂp��g��Ы�� ����@)">7*�2jE[p#�m���R�����|�J[��Hⓐ�φ�;J��4+��s5���$��]�R6���6�Q�t��b��#af�&�jT����TؑxБ$l�?��N-:��/DR.~�Pz2��?�o3�sxA�����]$Q�=�=CV�*�^Х6>��g��~���Yxı����֕~�\�j|��TU�0ڱÊ���W��$ץ��<8�{U+�M|B�� tk)�sR՚+&��q�Ā�%��>N�d�?���(�Ow�H5֐��?p����{�� �������H�f$X9��rŔeU;�F�V����:7Du�(�Y.�O(c��"��	uE��U���Ь���C��#���p�j��$. EJfXf�V�ƒ�7"�N����v��f�T�U1B�L�a�j!K�B�?����H���
L��zz�1z��-����RxĚ[�)�Yd��u���tA�����9���?�%HՋ�)���--����/ ����M�5�ˈ ��+*1��z�y9rjn�ů�x���O�]B�8?�J1��4�n£�o/�]G�������V���-� U"�Lx�0��i�~��$��� X��]�������[���l]XJ�����C�yF������a�=���0�����y�d-���(=b�)Ҡ�|�!�.��k�f�@��r.,P�:}��М��A��j���v�C��[Po�VL�	@l"2�i��B�������CK32�*u��vj���P�Qsm�0��uN���
�>q�x(��fx�-��Ui���n�4��!7��C�P�w ���00��^���h��Z4�~��KˇG�e�ݍ��	,�p�d�me�}�L�TՐ[���V��fR�r�� ��ʨ�c$��l�GE���+��]$!�*���I�a�z�a9����fP��68}���t�&�����`�5����N�
�G*P���#.E��L\�^\�ceY����j��!H�}j�+EO�@����ԧo�T=[���.�[A�JȢ�2[��@iL��� ��$㍖���S��يA�NA!ڪX�aW��-[:�\A`�H���O�=�2�c�����ȫ~���$�j��Z������Ws�"k~t�H����2��_N�ӖHE�e�ӝ��y�Aspt�uӵrI �AO����̔��Ͳ�6IN������8	�a�&��̍'1`�fL����L5�n>�x�تg�X�N���+^5Y�^$���8�(,����ID�l�V�s�����;�㒧t�j�G>DK�V�Q�|�d"X�1�"����On���I W]�PtÇ�/����cZ������I�H �|0[�PO
�C�Ċs����Z��-��`ٓ�K�� K�"�*I "�ɒ >��F��	}�в
�e�c~�[Э�X���I#�;nd?���_c�A����s[��g�*�ؑ��jg����ToP�|o���#���=�>��vN�T]'t�}���Ё�~�#��Cl�W"'_��<���E�e���J�+�]�W��q�N��ot�o�۳̍[�V:���pdxc%���ߙ�����˳��\ �_Xfd��W��kU:��7D���̗�������UƐ���k'�<��Z���1�M
���<=�@xu��|r݌lr�CX�8���m��j��F���B��q���1V�2�;�1�L�;<u�:���2���a��]a�}/GR�|6�_ �TӍ8�4A��L|��V��,�Y�h��R�BE!)��b�c�;���L�#��>ꋽ���F�:�Vw1,�;��TB��=� ��僝�`��_���hi�]�G/VhMZ�^̳���=���}�r��f�F -U&�\#�ð�ۤ����)���n8��f��J�,_����L�O<�z�G�0g��ǳ�f4� ��0jcG�-��1݉��,�ۊb����4'h�k8 "$P7����L����9�z�c��!ʡ/����@TT���P�|����+&�5���)�O����ے�'��s�qAL�1h�s�T����a��A������ kg��T��^z�oс�ۜ�[Φ��(���Fg�߹tA��� X�4���5�ŶFF�Y5�_"ܣYي�ׄ��'P:�!W!'�6�IFr�m�Fߓ����{;T%K����,|={�;�Xak�|�&��{��H�Mm�m&v�to3�]���m��g������{ arF!�`'�.��S�OdFf�ǖ��T!��� �-GW�@��P�քM�7?U��`�4#5��	���}J��'�֘R�-�Ng��>Gȥ3}�B�l����/�~F��ջ�����M���_���| m�h�����n���0G%	�]VG:E�#)�,(���P�= !�~T����b��׈�˺��|�
�+��H�0�z�Ԫ��t`�X�,�VAu�f��Z�DYG��T/�K�*k-\����+��'���86�� ��"8��(R=�O�FY�XnE��q�d�����Ȁ>�u!��Y��̖����)� a�<�m/s�֠M�\8�V�H�)lbV,�w�mޥ8�E~	qp��B�at���5�g��FO��I|��'��)bo*���*��бJ�>xCV�7i���`�tD��k�'���EF�'�%Q��܎�����Q4@���W�Y�F���Jkꈹ ��9KB_�9�tĵ<^g��I���b��	�yjȗ���� ;?u�nX)rA-���Q�¤��p��7��|'t�uH�wT���ZlW��`�t���/f�w.�N�Y��zDZ�h��󽲂SZ�Y�s���&��PO�k,,R�F5D*� ���_˥I)��G|=Ѿ���Y���E�x������Y��l��U���M�n����N���VLbRTǬڀ�Oe���e�3-I���N�8"�*Ydq3gge@e�P�/�έ��Y}�a: �l��䰢DN��;�Gcԓl��7�䷄U��v�� R�9��w�Gv�OTQ�W��ڙo�?ێ����.��0֝u�I��$����e���l���d�L�� �'��hW�/�OS.�|�f�P�!a�*���o1��Z������n"�+2�������Q��y��y������Ԗ���j�{�'�>C
h:�VL��Uc����ŒQz�ҏ�uv�Vjh�������.p?��)�9+񟕑�8�S�bf�o��ؓU��9D}civa�3k�fu�u���b2P��"@q��4�T���5��+����	�ܑ�mQ��+�'���[~quZE��ӯ�����6��5��'3M����2�,��{:�B�%73|�B�f��})	~���R^ԥ6qA���+S�j��48=dL�м�٥�%ԁq��~o����ϣ���e�sYi�<+��"L3�މ��V��\�6�O!��:�1z,�C��^fr@�L��
�I�
�v��wi�sI�o�*}���	Oz:+Ě�!@B�7T�C0����
j�Z�g<k�3����_�`I�4��Ɖd��WM�$A�!�ؙ�͌��%��a�0W�u]���v9�u>�Z�9�NV4��7�e$VV`\_~ShV�\m���������
��4�@w;hUq�,��rD���0��kcJ|�Y�����9�2���^Nn8d=�����S�j=J�}l�I�.m�A�tK.D���i�,?�w��e��.���ܤ6'�TW��,��F���Vڿv����+Q����;�W�[X޻"�}��ϙZɇ�y��)���XZ�z��e�]�э�g�&zŻ�������*u}��=��EȬ�_��Ie�h	i�p��C>�qr���X���+R�l۫!��c���7����ȴ����ȫp��!48r=:j�˲��`��*^����l)T������P!��v���I2���Ϫ��J0Mu3�E���� ��B7 � �`�Wcz�q��X�`����뭦�;���ű�G�ݘ�=`��#�k<�ywZ*�W��T*AA�z^�Z���SՑ>YN+�_`u�2O�U���Mj:RG�8vw�ҍ�S'��*�#�9<�~��Z��1�Dru����X���"4�pZ�(�b����؝~')��&�	���c<��\I�{el��	0z�!9W���$%+M鬋�l�$��!����8�A��gM��)>|�U
@�AQ(ǆowkz3�&�%R��B��d��:C��rO�$��{�5��P�J�\.��SW��%@�7;�y1�X��p�L6�23��9��_v��Į�8��&!>�B������Sǐ�|4;�%����s�:+`x��4��c@'�Vy�8;6�oq�n'��D���F�¹�^��(G���������0���1k�����������"���4&^_4 ��]�zu��A���@, ��h�����:�L�CF�E��uǳyQ���T��%\M�<S��Gv�
�8|�N�@���2H�PQ/*CD�Be��;DB��P�\�S�5��_K�)x|fR�� � 4*	�y��a*�ݏa#����A�i�>�g)�y����Z2���YϞ���[���>�X����X��0��wJt9[?�h������+�I�ʸ�-f�M@���ӱd�(�Iڹ��F�H��.\���)I���)'9s���o\��f�B���Ѧ/}}�tH#��=8���tV�	3�mњ�	�
�+}���3!�$0��i�°Z�����Pߏ�G[%Ȋܕ8x$�U�N��g֪�H��smS'�J ��[�{Λ=�V��q/-�fI������wѱ�vW��8�1H�����B�z$3��E�y��5���W����w1� �tw����'#a���ﾷ=�ֹI�=���t����ꮄ�^�V_�cs��؄��0}����RZ�v|}�$�
;$R]�f�Y�J϶݃�Gʆ�y��L�����GRm,=$^c\cy�4��fY�$)�g��M�岚=�0Rk��O��#���+�dg�/�iX�y��-Ƥ�U�V�
vڴ!���I�N1�ч��퇰 "6�i*�0��TG��!�C���#���{�WxGmp	���;I�Ρ�AL�M����
����^`.N0���)�l����o��|Y^tq�9`���$�E('�&�좤@4����o��C��7�b�g�>v%�ޭ�rH�#L��Y+�t|N[�>WU�=�´f��,��S���&n�7t��o�5��c ܫ~�7�/C?�S���(���H�ܴ�G���M4�O�Uoʹ|��fdv�`l����c=F ե��F�z��B�mf���LiK=i�t�g�-e�M���Y(E��[��n|���0i�N$���n�\xWc��H?�5��G�.P;��-�W�!Y�����t+y���l�ê�=�O|*-�LaR��b�k�CTS�3�I���$�`8l���\��sG�d���ќ빿g�l o��FR��I�!�6f]}
��