XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��T���8���~w"��iS%�;	�>w�G$�ŕ�X�ޯ9�l�ͱ*��Y�]_A�s/���`�<�_�������肄9�F�3�/!$�fԆpk��i�cL��X4E7�G�S	�?�ꮠ��!dx[c`5�{-ב�^x�O�Ǔ�l��Ý T:��+�7�O^�����*%"��3�G���A�B�?����!��>"��⎾��� �׌�E�<s$���p�^�vNb[��{}0���H"�0
�e�Axvƛ��fg�rO?���|:pК����I��u[N*�ɺ�1H�tU*������/�ӝ�`�EJD���ݓ�&X�̂ќTJ RH�0��CGf����|^O��F�&fO����F�R��I�6m�U�����/�J^��_xADD �Yg�\#���������r��Z��廊�8e|vX�J��ytI���_4\-E��,I�x�����J��r߻��,�-w�zw���� Fl��Рl���Dc��uA2��փ�O�+Lz"��{�(}�v�Y8�ק�7���@#�c��?>W��K��XZ���Vi�(��ث��>%۹��$�0��I�|}��:���t�d(*{:�h��A�X$��?��b��P�Cq�R�9�(���å�/��48�/w��ƪ���G>�o�ݬ�2K ����?8����Zf���M
3���q;U8ҋ��������#pO��?Rh�����2)(�l� �]��9JW��}�l�q��XlxVHYEB    3c92     900��2P��o��S�cWc�OJ�����C1=�\|4����rhv�\��R]��^�S�3s_co�5�	��S ��3˛0�.���R�.��)/�P���v�\�<:�v������;���Of�����L3�H$2�G�p	�r����!'y�"�ִ�b��s{j[k6�̂gb�HH�X�Hqv�f��Q��y��z[�Ƒ��NUx� ��%�J
9\̕'8�S��|b1;�8�u��/3���E��x�ot���S��L��'F؏S���`7'~�߁����yN1�P�����8�:����A�ލ��5e=��P�g���@��1�v���շ.V��#.�,���Ɣk�gT�j�����&�v11�x+�]m��و���$(@����i��b���TƮW`?�k>i��x6D�9a �W�>9���~Bg��f�t�`i�w�I�E�Gĭ��͞�#�h�>U��N�u�o�x���e�6��O<��l��Zya�H�e�&TM�XUqJoN�^���њ�Fھ������3au��x�5�]�h���������J�<O���̯Vr=[���=�g0q����]���M�g@��Y�vR9��6di�d��ӟ��Ϸ�OR���U���mhtb�N�,4�.��!�Zu��"�}=vJ��1p�s+
@S� �o����C��R�Tybȿ���Z;��=�7q8\�ˀ�,������j��@r�@��5=�:QhM�2Nm�ؙ����	��kͺٻ�;�աz�V����ܖ����ؿ��YL����$M�i��V�����k~m��HIs���2�]�m���A�/ʯ5�n8�E�Ѡ	�
�7"��R��s�sF~E�����u�pƬ =���\l����L����M���)+�\�(��{׀�2�<��ȔF?����[�37X2���nYed���/�����
`�3e-*���H��u��"L����v@VA7�T��Z��R����R�� F�"�
�fn�Z6���a�{���NE:q͇n���L^%�ViƏڵk���T�h��-�5IX��dA��O���*q7�0�c���B��L$v/5зZ%�js�c��ۙf�ߛ�0�}����8���%`�ţ��gC0#[b�;pQ�� �ˆM��e*�#���jƕ�p��왁y�,X�$K=%v9 4B{��Q�;މ)����/�}ͬ�"��}�>��o~�ϊ��M�=ǉ��E��Њ����� �t1~��h<k�A��'�HY�rDs����2�_o�g��kj��.�B�ƳN2��i�H՜=���b±��1�q���0���Ͽ���{g���L�4�T���6X��gD�Ӯ���P�/���<��m�N[����>��F���v�`f���d�l^^.�����#@���bL׹O�64��H����pW�y��E���eF��L§9epmk���i�z�#�2Y�W�q��J�[:���dEַR��=Hb�y��	�7y�Kܻ��g8�^���my�(��wl�38Kǻ�]��}.��넉�6)��rf.)����g��2�ec���V��jI`�+�Bm�)X��'���rCs��^���7&�Y\���>F9\S�cN01�OS��3�r��+��v��=��@����Y�?o;�
#�ID�w����Y�fKy���Q�5[Q9��(`?���x5��Gh͍�e�]��[tJ��r��̌7Ή�z�����~�z��<M��k� A�9}�4.�������?�DW��FE(huߠ�[�Ocȿ;9�ƹ��³}���|P!�.��?Bw�3�d�S�e>��2�'c�Qc��!d��~qn;_?=���?{)�fi��O��=�Jc��3�(�\�ޞ�c33}!�)L��8���6�+�B�/�"�R`�"l2��s�E".����=�	��-��oL��ʢƓ���U}Xh���J� ��\�{N���O����x��.S��l�^��tv��g�N}IӓS����uFc#˭3Hr ���M��0|�d���8�����\��>d��W�D��Lg�.��e����h�/�����(�-;�,�~Aش�� >�� ��)��&��;Q
�:g�̆7��xO�]E��h��}���v|�`��dh.ŭ���2}��j_��2�<$�[YD�Q���X9\>+�Z'*%�a�;����b�����'�%�m�rfD�|c��ٓ��D;܏�U�}Һ��)�4����K'�6~z�O�h b