XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��������*4��S�f��~����	{k��Q���:��P�?�7Q� �7�)���wΦ����p��|V���	��.<��)��0�ɬ�y�J-q:=9�A�-p6+�~��5*a� M�}8�Fp�\�E$�y�-#��d�05|�t�P�PN%���s�9Nj��8�pk��d~�"�E����U��^g� �O:�����Լ�-.�.!Ũ��ն-��;I@I"!� ���� �Vq7v��b0n���.��p-�;/��ʫCq�f��"z�E,���!=GDB����A��s.ev��ﭧ�Xӫ�0���|Â�������U%�'�����۽G�u��k5�֏�2+����9�d��b�u�Q��)ǫ/��MF|�nÀ
ry�|��@��xR�i���i�X�����h�sKV���1������R����KG8!�!W)a���g	��0��~�2�H�w��PQ~A�Я����?pj/�"�/^��4��K��ӕ�T�!V{����h(����[���_��En�E)s�!_�:��H �Ve}<����[�"������������-���!�&ӏCJ�/�R�"K�	���Ih҂�����o�^��G�
k;f��)h.%'��<��%��*�Z͕/�eVY�m���=r��wX}cF!��,�hX5�Ǿ��#� ^��Nx�m2������49�������^�/x�X�����u�ҿE��!�'��R�)�q�)�^y���XlxVHYEB     9cb     230�Rܕ�F�t�C0�G�"0�7��>"��GL�N��d<$ ��Q������_���]��zSC��roMFV��eP{��\��i��&����^.6[��`�F���;�� ���CYnf�A��[�1�Ԩe!�'H�WvB�r�觖�^�GbI��d.Y��"S����F[9�Tւ��_�3�o�l߮ނ�%ٌ����R�kys�:�:+Y��j�}�خ�yε��CQ1Y��ǥ�T��:nV�І]3�jdc���L�l��8v��g�qM_N@;8<y�n4ͫ�@�.��L����E��=�ɍ��3�l���H�1�L��MO:?U��s��O`��JP"�Y�'7J��?,i��T����^���.�ʹ��a1�;ZT�L�K{��\'ﺆm φs��epˮ#�H�\���M�~ϴ��p:�ؗO���6KV�Nx��wx��c�Y1�G�2�?�����De�%+�O�G�Д!�w�)���Ez��('3�Mx�D���]F��-e�������HF��������l�1�� 1!]*:�}�<����̈P�Ie���w?�