XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��4�ږ�}���E�j�xl�sՙ��1��g�R�τ�$D�)���շ���p[� r�ߝa5��!���|woJ��x���>TL.�����<���4/���H�!޶����#U��$W����3�U�_-B�~)ʧӱ�Y[�u��g�D���%�El��E�������x�}t���G�S}K���9�.��i��a>��h-��NkT��n?" �,�S���ϠPs�d4�Kqng�ؾ�Q¿>����{�41���.��3�:DX�SW�ݲ�r@����؜��L�3�^�|�{=�9�l�OK5�:���湗y�`���q�_�c������-���~Ps�1ֲY�W\:��Dv����4�&�u��Y�]��4���d����kP��`;齃,�l�����j�>����Ǚ`9c�,��a./�vy�ݴ
%CV��#��P��l�lE�V�x�<��L�)��V�0­��
�1pv�`��p��r�x$Qh�|~3��M��g�Ϲ �0��ұ�Ʈ��0�`'����y�dг_*�և�/�A�-��f�#��1���v�����ǚ1�7^2�Pe��1�Їn�^6�s��~��<�C�%�)����:1%F'Gx���|vY���Yc˩�̹\���my�cW@ ��Y����Nk�XU܈��$!Е�I��E%g��(��n�7N!�v؁W��Y��k��<�Za�([H�( �dJN9^��$c�Ϳvl|J�v��qTd]�@�.A
�� ��XlxVHYEB    1569     590�6,V����h����s��:��Je]�Q'�jB�*4%���9� J��I�j�o�r�>[Pg|H8�;��Y��2�W����Vc����	(ƈ!X\��G�C�E!/FN�_��E>L.0:_����DkRl<�FZ�|t���]RFx�N�&���;.��}C��&���9�k]i��� fDX�T9lwA�B�&�F�Q�D�'t�{�����Lk���Z&�n����x��[�,���s�����('��X�TQ������f�c���ז��D�'�.�Ms��� x�<lZݓ2�Q���f?͂o���ȫ��`ixN����&��Q:i_x��?`���7Fy|~1�����B{e����ل��N%�sa�����$��<(Հi
=��c����u�Tw5x������M�ҽ-IՊn�7+����pZR.$��	�<![Ϗ�]�cr$��`��w�~un�IBT��μ��'�N�ֽ�� ��n9p\�rD|�I�U�����y�Ђ7AEf�.D�rN������+�Rn7U/���u`��ٸx�^�9����fʝw�J8wI谱'�����@�H����s��}rc���!�E�cEѮ�o�̔�����(��Y�6����2�:ݤ�r`;��~�LB%�n˫w	����
��%w�8
]�����E�����'�N�빼�pNJ���\M�V��9|Ti��0[քkB6�N!�A_�	g.�l�x���([jJ��_�Ny�''����!�؁7�R�
譿�d���y~���7� ����nq�<�^`u���00#��s9U�����S���^��7r�!8Y?�G����Hkﺣ����0X���kwn�=J�n�H�� O���LRH�'�1�P� ��c�9�'�i� c�,jQ�Z�2��&9,�Q����	���0�w�s
�N�Ⴚe�t4G���Fv>AĘ����*�D:+����$`P)F=:�ڰ����2�3��|�/j@s�[i��>����b���� B�<�!x�bl�9x��IzћTلC���KgH�o��N���07�;�6Y�C��)��H�R���_��SAṵ/b!�8�:Ü�4U��rlJ�[G}Ѭ!Kw�1��^^��טqn�����"\;0<��S��0�jݴ�:�g���Iq>���mD+@��IQ�������L��~��$ٸ䀭�n���c>^3sP	����=b@=Ј\��ݞ�"6�ބ�Z�{�~��,�JY���=Il^��F���_ޝ9U��t@D�)�k�w�"lDdD7Tu�����tA�^\X�����|�<��3j-�t�ös�1/��>���g��j���\+�"�k�q���z���ߩ�]�~�