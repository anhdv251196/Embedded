XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Q�>G����&� '�<+�sn��T/x/��*�
�4a���d,rNB�����=�ȐL&��=c����(-�u���GB@��v�}�z��ľ���"ʏ5����+	d����1I�,�Zy7��T#�gR��[�`~mN �e;��jJ��bX�}�;r�Y�Ǫ��`�v^� 9Rlɝa����M�c��/p`��׆�X���ٸ��_9�7�����_7X7�<�ӟ���e��x�`�lʗ3U������qt�L��Wq3JZ�kN��.�f谒����|����ad][�����vzl��g@�=J�N�ߙ���*�12�ц�-�hzHi�/���=���V*3��^�o�Sz��rd�7XbQ=���m��"�g�@:���js�AaJ��pQ~;�GN�%&9ژ&�jnt����ϋ����F�#8'c��D6�s�rk�<�+=��w�7I��f��e���hL�����]���c�G3mޮ���i6*�#�@B������?�G_�|^en
Q�+r2�E!�Ӊ�O� k�\}8*��|i��-�ʜ��uw�9~m:��ֳ)i�&�\�>�+B�~��0?�д��݃�fDz���v��|62�e��|�ʾm�0Y>�n�xi	��,/m�,iJ]��v�����f�j/8�X�2�I,_4AF���$��[�1O�e�kLpVg�\�g�(�՛�(������H,�[�W/KW���~TW'&q¨[^����,�7��T9�&rtn��XlxVHYEB    1001     490�(�z���V���o�γar,�0���"���"e��"]f�dP� �渦�9�fB=_�5z�g=�=�^�F�<Ħ��-"h�j���3����rblr�*�_�dj�4���Z�������|��^�vGr����\ء��gV�G�� ��!;x6�]Ck�k,��w�!jxf.��V ����=�tF�jC����֑B@�Q7����.���C�])>O���\�0s����q����a�t��a�
��d:�b�3�KE�x�#
`5����7`e;&�q �_K�������.�m[����&I�U��JTDeD��0G�H�L'�|�&�Q/��䡾9�Í2��e&1�2�:���msȐ>X�XX@��o�]:�D�q?/��Od�@�'D$ƄGa7횵�]N}�����cM+��N�DS���2��t����W���`]f	�2��+�WDG�@�Լ�O�����J���f�䌝߈�뙮`�[�Q�{�:R ��r�t<,*���fk����oAD;�t�q�q�a��!	JV��
����}֬:���F�:�A���Z�EsF�5�����۔h�B��O�N�:* �s�2�њ1�v����+�-�B�ui��^���:M�d
�r	����h\�W�S1�<�%�O�l�� �{��M*h#���q��f����y�q�أş�������H/��0Y� &���`��������W�
������%�\����_�z���pbF"栋H�zd�0� BB��i�ٹmr�=�P(������rrh)O�X-��	��m9g&�W�)�o�J=J�$ e9k��r����끂�*����ih��Wf<1���	�S�"�5���"�V�O�ǣ%B�Zk�S��K#�#`C�� �;A���Y�9��Fi� �g���IK���Y+�~ՙ^nhn����C����>!�����L`������砈�����h�8��h��3Q���	7�{�U��B$���2j�|r��E���]*{�u�_���k��%�-Ϫ��F���^�"/�-pם��=�=q���KC��dl�;E�1��ʟ�.|�>?�%�m�BFW%f(�)A��	/<�jĚ��І����$v���|���Ч�x���d�� �