XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��u�֊f�b*v�"�F��1��Vzd��0lJ/'����gTH 7z�G݀������5�"'��crb<��o�����5�3����:S���t���'�l&��|��X��Z�ک�L��M��2�c!�����Jn��Qѱ�S�*׀|�;^c�4K<��{Vx�����H#����P�*,a��ò�%���x��Mu[���5n�u��I��P��z=L`���b��N�;ǽ��+g!�r4��I�$jF�����ؠ] �۲kp���e��j��;��zn#����# ��v���}��	��B��B��K�J�_��^b�QcN��Z0����1���|֏B1����HC8���穚>MJ��3���qV�JDl�c�wڠj��e����&���?F��ē)v�	�H�l!7� P]nUW�u��ܵ#�i
ӫ<���L���=�i"��7t'�(���j�&g��Z?l������m�]5��0��F�,��F2���T��g��r�b[*��۱�v��}�'ROno��<�L�uWn93������h� ~�t���߼����V	~�r4���w�,�V�1ez�?�sǋ[}�����I�X�Gyck��9��_.Kܙ�C��<���d"��DYے/Ց^h ]_A�v�1<��ݙ\L���%�e�;���amχ��d Y�|%��L�"�j�amW�����R��-ߔ.�1E� �w��"sae`��*
VY��n(�#n[�S������\?.^s�Q���έQE*��+�L\�X]XlxVHYEB     a7c     440S�W��ύ�f�CU6�l����+��&e.ڹ�J�xʄ�(2yY��.}M�����0�s�@�b���jدӒ�T�m@�3��Vw�O�*�=�K9+�!�/F+�Vϧp.=�17]��'�P{��?�ri�Tm=��(r2^JϪ��_ˍ���k��5��8rll�Wk�x{݊$�y��8�WKc�P�]ZZg%W��W������Zd��JK�e �
�RN�4�-�zL���� TѨ�����i1�ʦ%v8���YD���S������V�y	A�Ρ2�<�%��4��ц�E���F�l�oH ��[�S�ɤ�=�l�_����e ����;JM�\r6�R2�/�FLh�|�;�Ӛ�p��5Q߁N	I��o]ă,�ƻ��{+<[�񖾾>1�����ObG]����'D�L��{�Ii�w��L���]Sz��� �M�&Rx-�
W�;��<}��=��8��ؖ;̯o^*N]7X�B;+��~Z1;:��8j������F�m�K�u����9�c�K�B[K�����1\������6C�?���=g6������0���w��T�|,����5:�O����ג�^�Nϒ)vJ�825�y=�Q�EP�&0տ!n��>�㽻�,�W���3-w6M����%Yk.�B��ys^�GT	)�Q���Ri���H6�n�"QR{'.�r�+�hm�n#O>}-��mHuОpA�ti�s����Y�kpr)���x���_Ɖ��C`}3>KN�n;��r{�	Y�Ve�a��L�J"�֏o�b�h���5�z��v~���F��ݪ��@~�6�����7�2Z�"o�#���&���Mn�I ���C�p�<L>�\��ek�
#������?!@W0�7^�1�;
y��%�8��h�P���F�)�f�~w@7''��f'5c5d���y���܍��
����P"���xq��M�§驂o��TZ�m����� ��Ȁ7+��cx�w0�	�e�������}Y�,$����cx��$t��(�\���\��o�憺c�4se���L��o �>*�H�