XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���?��Mg���2��Q����t� �Iъ츷*�^�@�z��T��4����))�`��\h6e�Wx!SUL���hSf���a������y<<JC���+�Bz,P���Q�qwS��*��o�P�&�h������^FK�4�s�Fp��w�NW�!�@��g���&�x����L�{��H��E�0����v�Oc�'ɑXk1��&Ǘ����L����V?�����;�;���F��,�h�Y�ZV��t�[*�����Y�]_��p�Uc����Q��h�ɼN���3Q��S�z�j�Zz�AD����9(�A�,�:�u>o|�bm�K�8*��u;�<h�Q�z��tO�r�=����[�=H�}-���~"��q�9���G�P݉��/��p_�Q6�:���}�=4Y��5IV��7�N�e�6^�����$rC�nL�h� �����	�������H���/HTԛ��R��,P�ײC��	���/NƱ�Mv�"�X�▒��IX&}ep�_6"�2fѾEѴu#�5f����I��B���5j����f��3U9�r��{r\u)������t�>Q�m�)��r���Q� __)�@W�kN��n87/��S2ށm���r!0� ��P���N|��k��D]�i(�8v�~��$�T��k�F�M��al�R%���u��+)�|E_I��X�|��8�w��9��mϤ��07�%�Y���,�#���v�j���AIQ����4�Xe�+CX�Olf�XlxVHYEB    41c2     c40����×�;c���Y��5���D����¹F�J�5�h}�"�G!�6�9F�����՘�˔��g>
�e�Nm�]뚽��=�>8��Y=��+?�o�hvx��=��t�)���?p�,�t��1H,�:�����'�^]&��S�8�@E}�/�@_�+�ӄ:]���1ˬ�]5��z
��ҩ|��ϧ��> ��q�7Y8�ZA^���{��T>e��]�2�P#�f��]�����*�N��������
~�+f��I(xCZL��`ٗ掹d� ��s�S��M/��[�VܦY�U���WG�AEPR$��}+���� �[O���x�)
�#d�=�E�V������s�:���I�7�_�~�c�<w�;��ۧ<p�Z%)
��D}OE�v���
k�lonz��_d�}E	�����JP������:Sy_�M�Lk+ +`��p�_��{��;��t���ꦌ|@z2]���_�	:�X�k����j�C	��_s�v���bc{S
ȣyd�?[�����98�%qDv�I�c���7�`�E.�2LT�[]];ρC���ך"�(j-���9��_9 ���i]I(���,1��Z�I��R����� ݡ������q�%��U��Dу�=3�K�=$���iD�y�e4�r�k�q,���]�嚹ԏ����l$���/&��}jK��y��x9�ҷ�m;$HB�v����D�U��W�M���=�XC���bGʮ=��s`付Ύ�X�TQ�*�@��-�m��r/�b\�&���i�'�?`���o�Y���Y���=��s���&�[�yy�d/�����]��]#2����1�`_3L�[  �2���M������\��`z��W���V��1+Vx������038��^!��5�I.������$q���\�u6��dƘ�tׯ^T�Y�����5�1�t�ؼ˒�����5ߗp��Pj��;]g�4��eS{'3�H�>q�;ZR�6�:�GCt�k猜H���pH���P��:�^��0ge�8N%oy-H�!��Y68������!�EQ8��D����9���@�#���a����XH�{+5>��m�N5Ԉ�~��o�ԧF�\8f��4;|���@�����`JWoL���r���ȿ8�&(���O��6��)|���J���#6�=��z��-�~g��[j��*6����'//P��>mV�#+��Iw��й#�N1��V� ���x9�È���
����j����%�e�k5��_տ5�'�����A{�e*{pTL@}���3����t����!^��,;Hj�����6P�y��s,�M��R��J��,Q>�DtwQF,���V�1�r��4���5��H��)m����uj��Ș�P/#w�YZ�j#Z���fG
cI� X�I�2�D4dL{,jJ�?6���6(I����<�P ���_f6>��D�@�~�QU@ySC[��ߪ�ř������+{��'U#
���:�6FZ�����
y��s�y��4T�Z���Z�"7�M �i�g��ǿ�b�%�9�,����%9i��rG�]��3��bB����nH���1�7ɪ���i�\G���Iܔ}cp{X�:0O���f��B����Y�H&���`tu{N�kU�z�bԪ�ø��f]z�}i8��Hq=�-�a=7���
g�QPc���Or�����S�К�%&wن�/��$����.�'Ƿaո&V$M.u
���Q�;��M��n���H�ˤ�{9�: �� ��K��=f!��RK�؊C�ܹ���l�K1�v畴�H.Θ�2�C����@/�����W=kN�+��*l��P�#v��o
��}�mTK� ��`f[]�Z>�5��:��,˶�|�깏��+�th#�4\�	�ۄ�*aqlގ��=�]��!maN��u�+�r�U�5�>�ˇ���N �M�"�!��m��Q��b��$��+�^��S��bW�C2�8wQ��췙PQ/���Va�R|���Lǡ[�P�l�x�5�қ�at� ��o�Hj��}i��R�S<��K�/�[��E�-h�>Ƴ��E���"�8	�SԂe�i���Nej� X'�yL�`ʿ��������>������ӉѾߟ�`����k��7;�A�V;��o��q��R�Fn���rԲKY�ȳr�� �Wr�c���^�v$^��A�d�(!7���9�������R�;�RDL��R֞x�Ƥ��-��7X��01�Ӏ��ӯ��� ~O51m�໔'@���Z9� ��q��DN�`I�m�M��Xsr�!V�@�V�/'\i�Z�
x]�4�&é��"Q �p���6�l�(S��*/0VN�	J���q�җ2�����/��O�C�Ky�uTH��WfU�D��{m��y�C�,�������3�i�Y=�o�<|c�6u�;*�������E,�`B��atx��3�4���.��%G�?QČ� @
x7�`&Ua�I�6n�'^1?ONAr�K��c�LDIMi�?d mȩ,��a��G��\�����s���&1��t�d��>q�r�	YNxk�~sa�������gb�'ٸyj�Oy�7.�1�O*�}E���䰏��=�����\pZ�;��,���2 �����$�������X�볿by?尛��s�0�H]گg����ΐ$�#�և��׸��w�����S��)��G�6FK��J�}� .D��\��ƹ��f��Ώ�+���j;.r*!������h�d�}e�lc�bt�����%���P��^�=�\;� a�Z�¶�b����T��W���g�
k��A����Qf�҆�	Ώ�L(ch �����DB�U�g߃-�� W���_s��a��#�,K��	����:N~�<�<�H�J��B�2�d2����jt�U�LV���QS��g-����s�A;F�ڎ &;�u��}�m/7�1AT�ۡ��C�@Am=K�Q�!��S�9��y�$.=ZJ�:ئ�}.K,�8;<�"x������jJ�b4�x,H}UV��>��ﾑw6�o����H�^)��>-5G