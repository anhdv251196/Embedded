XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����`��H�whu �
��9��G�Xbe�YU�f~	���^-�/3O-�E:��L婉|�8;�)NyF�ģ*���D���]������00tXZW���I&�`����u!� !`7Ыy��^s���6f|��g? ���,M��WVj^o�*t6JڂO���]�Vy��V*.�xeg��V����TW��)�������6�=�M�L�x��	(͓����2'�d�颠���[��)�X[/��-���J�O� ��x�7��ab�V��0`r#P�slY�oQ�s,�=�e`�,7��m�ԑ��� ZIt�b�n�k��@/��|�'6D]N9(���n��2�6;>z�UT�U	��u�j_���A˙�Egث��7��+�x�=���m�f1��e��)�	(k��F%�����T�q�o˱Lw�|8�k/T۝��[H'���s���m�e~FK�,��ӌ�z�Z����+���e�^gTj�d�
�}1�i�k	�4�"�8�E�18�;�j��?�Af��/c:y8�Ew����|��X]e���3�H.fh�$��F{�Ӿ=\���楜��A����u����BD%:eyq_3��W�b��Q�4
o=xz�bg�U1����h����x���]-�N/E�q}�M�>2WR�����(�?��U=9�s	�%��]���E y�sq��,�8c\�z�9+�x(��P�f�Ê͈�[沠 7�	sM%N���5ؾ�+l. ��~c�E��At>eq~�B�m��i���z�����XlxVHYEB    3541     ca0���6��i(S�OcI���ހJ��0w��5��ݽ�X4��l�3�\;��3��>��6���|��	��m�F(���1��+X�D7؄��0�O��3���k���lJt�dex��Agg�E��V��-��Q��-�c��I�2^xLH��č�N�cA��ߥ�&;��c/9����s��q�5c��i�zޥ�V�ן��N�g*$T���g9�;Mp]�ܐjD�����A.;�k}�vo
~L�6�M���uk\XNMC�&�K,46�a�EK^E��(�Q3n@�����Zs�G�lW��W!Ɏt����'u9y�];4&�G���o=%7�`�Z�$����2+��3�k�<�H�ڸ$�M��Y�t�̴.aصw{<Pm
(�}����=��%�����IV1�J��"�O�;m�#7V����O�Ƶ���͸�V�1�u�Ԯc���2O�,oi�~�������9}���Z�У<�M�h��o�(w ��S�m��M��\r��Q���5#�37�΢�d��2��V�ׁ)�����s74Z��C���6u��&tD���{��R �_B�z?�[U����<J��,^��7w�|��	�['�^	m̣����+YBt��[n/�NYF��c��G�z<�k����7�qn0+�V.��#i�DAgӔ�[ln���r�q.؜]���@�)q�rB;.mc�;e{%��ǹ�6���:�h�Ғ렳I�Q@��Κ�

���t�'�N�i�O|Bڹ ���2�)6���Bm����䡽�ʍ����iYGh�}�;��[˒���}�����M2'��ĤK�vځIS��PwݡWԏ�++�R�~��7�lNH���\(��52�M5
;XV�����v����$H8��\�T��^�r��)0bY�V߯v������Q�������<���Z%c��w��a�1���S��~IW��VUi�73Wx㯆/ݬ�(�qF�q3��Wlzyā�Mlj`^cHb8gp5V�G�?��j���9�5�lJ�t
B%���]͏��L���z���H�^pC˻��m�lPT���:y�o�,�����HLwZd�f�L�32:�#!�NQּB�ܧ4�Ǆ?�aÖH�ȐQW��Nݣ�(���n�8���;�Mv� g������d���
�R���u&��{̓XN���֥8����������^d�P6#bd����yh_)R�HG��}J��,��r!��ǠKaӁ@�J=�uB�l,��D��*���� �@�����u;&�ϩ��s>`��4c�_�2�1Em;$^�IQ�����⎶F^�04T
^l��֑��0�����"�1U��6�6�<�u��올
R+�ORy���J��mkτ�
(�
�r/%K�����{q4z1��ʃ/y�"���C�P�)���.�:�!�)��$�S�BB�B�Z�A��=�Ӆ�W�,��h���H�fhG��j�/$�Z�W�E:+m��&�L���)����#!�1.S_�Q�e�u��;tNcP=ݜE^����EV+<�EԺ�@.V��Y��nG�!o:����S�Y�;�D�m����Z���:Q�I�<��P$b#r�Ux�~�����⫑Kt��7�ҫ�I �l��RmO��`�<���Au�lْ'�&��zNL�i�k��,������A����,e鯛�A[�Hn��0dN�mZ���P��#S�a&x�b�k&�J$]I�y�w���擫��O�a��!lr��18�6�4W3Y̦��x��q�) �ͯ�^����*�3Zw���3����Ⱦ����_��p�Q_ [��:�;׈O~=xԵΤ3�e�q�\��빪=�oy�ɒ���x�|r]c�Ȋ$=��NG�8
&v�7��V^�(91}ye&*H�;`Bd?'7�,������>Kt����y������5�2��S��67y��Q��L5���K�]�[����=#��	�r[/�k��`�:T�붎&��	)x�Dd0<6�]�����9��Y��P�R�!�r��d��δ�^�t}@�T<Hv
�]��iZ��S�$<���m��3M"�:
������D[��X_e�(����:R|5Wn�`F�<����e��"A�����yF=�t
i@ʔ���&A���'�X�}@���3�+�*A��]���v3��?~sf���U��o�o��G�.d Ux���;fo�]�BЈ"`�§���(�`V(x��v��p���:yH}�MMXF�F7�����i�1��F�����Դ�J�@X|�k�3f���đtA��������'*'*I9Q	�u��XƢߵ��4��%�����#�9>���s��-u�Ҹ��~���&$&�Auy2fe�*KQT�p��:���).X!�g��/?V�����)V5�������OI���M�b������Ig�Q5����W.�\����A0Ҭ�m�>HY"�T�;�It�F��G�����斯ݟ��,���c��qW����,$���x��P���Ǆ��Z��� ���`�$�M�R?%[�h{���ae�x]`�	X��Gpz���R�_��n���yn�|L4�����1�X��,�����u�65a�K`�͔�`�xK���a�d6"�5�	�&}����&	�R�eU#j~��
��?w�.�YH�
p����iU�&Ko���Dx:��0&-��m���4�)��g5��B�5�tPv�?�Q1�����m4�����$�6+Z{o8a3Fs+	�"@gz%���k]���[L�
��"z��ږ�THr��¹��q�+0��2���S4�#���uh��99Қ�S�W��$<�j7a�|r�fG�9bO0�WR.LJ��Om/�%<�H�l���ɡ�3 (������&V�e�����٩V���Cr$����'V�b7x㟢�:BJE�~źPW.���~����w�G�7VhI�x_��C=
5�*+h�x�+��H6��uV�EH[�tQ����(?2���&'����J��7�B
Jbe�:C����$g5]��� ��f�_Xt������;RI���]�!e���,�;�������*!�\�~�Y��Ex��V,C�D��Z��#1b�
vi
�U��H���jE����6{
ԧ��L�b1Fd��A�=��܁���