XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��`T���L���:�O�D6T�>�3�����^� ����&�
z M���$w�������j�M`�����Sg���cӒ?�:2N藬�7���*���:vkѥ��b�j� P�x�U���ds��^i�Ԯj��/l�!��O>�k=��Đ~��6���	�Z�_�C�#-W$��W�.`.X�`����_�M'°*ȴ$���+��v22��{ҋ���{�h�$����v�QEw%V�ѵ�t��t��N�����P�̽�	�p�Y�����Ͽ�^(d�]�|�ý��g� ��^R��ǈ�bf��g����Ch��s&�`��O8��
Z ����$���x�X7^�Uv���օ�Z�G;�q�'SUR{a�+E��N��O������[�J��8�S��R`�]�Dz�P�^oeZ�|h�`>�A�ƍ����o��&���M�7ΜeߚGך��zܙ��C�Se��=�$O��Y3u�<N��a�%��in�'��C�3l���yf��X��яyR��{�b��<[�A %�t�	�8��JQ�!7c��&����XE�T=O��ݮ�+xR�v� l'eS�yS���Q�1�I;ph�)}�J�m��p�ӯ�k0$�jt:�~� �W�4��\���I�g�d|{������~����"���p�$�4ac5B�g��������Q_ɽr���]����c�T5����^�����e	�#��Е�p���	���Er^�A�%m(myH�#+�uXlxVHYEB    5ff4    1040Ϗ�Z��g��u-.v�1e�c͹_
��-��A{���S=/녗hWt���8 �鏩M9�g��-����tU���x����u���{�4r�5�_͎�%@�!��U'�I��)Y"�m%�%��iVD�h?jY˸�K`&}�������ʀ�V��Ll�.������� ��z��CeyZǁh�ޒ�����{ `�j��E"����:��1AP��Fy��7��3���wo�D�ߞq�!.�!~ ��.Tr�9H�=Y��M�_��Ϭ����I+�����4�ޗ���bC�x�c�0X Q����ا�s��4�qN����v��K(Y�(}-���lM�N�NS�
��f����?1�����G�uؤ�M66r�����O���.q��)`��W�H '��g{fv-yz�{-N�n���j����W�p+:��dz�"|��z�Y����j�R���kr�y�K$�Dw�I_�[ԫ�V, �9�#�6G�u��B�]��Hq湃T&�e%/�9+yBz����q���p�V�li�Qm"��q��%u��y�.�<!�s�K�ľp��F7t��u;�j(�a�AnV�� -Z7�E��p�+�W�������9>�����s嫯�����'�WM(�ùo�s�V	3^�'�nO���[t}L$9�1V��4�m4o䨞Ņ:��C�Pxd�cRa���H,F���#G`N<�ƽ���Z�z���4xE��ۑ)�A�6Y��|�����`gw��X��C�狥k=����j�����1�CJ�x��eߌ�ν݈�oRU�0{C��2�a`s��{;y/��)��]�����44�
콎_Y8%a	eK؈�)F��\�XUd�N:����
���ǎ���Ғ�$��:���M��L���k��L,X��l[X��:"��>�=l��.n%7�&�M�'����-j����趚��L���%M��6����DE'G�ǖ'�`N�ż3"]stL��:ڤ!�Ğ���c8G�%'H|�7��YɫR��U�*�Z0i	�ӫ�^2[>�5p�x���߭:�/�+�a��=I����q���'ʴ\���!y�f�������C���x�>��ܗl�ٽ{��P�tVu��|�~6h��}N��.T���T��q貝����%�Cd�����9�����3�>\늋WC��Ǘ�m���I�f�ecO0��)�fS�ήTjo��//^�g8�sCTu��]��G��b��*�������I!v�"����,���i�F���h���!\Mg3�u~ŋL���.�����ͺ�߶z����=���1S�p���5AB���'�h~;������;\�fJ(��*����7��>��:7�M��<�U����@�����
�V�h&mzkC:�pI@{�M"^N��ü���-J���~���k5E������E@��o�U�w�b���J���	j�4Ԅb��I����P�x��p�`���H�=��侘Q���B#�J㣢S?ϝ|�����$��L`ėd`x0{�+�z������e��kq�X��8���T����K�V��x��1_0�y�h�n<[�/k*��1��RZd�,�4���>�M�=Ѓ�6E@�2q9��q^O��ۍز�o�C�h��X�'�/�B��@G
v�3�qd�z�I��A_#�q�+�G��ee���In"�6[L�׸�-��*D�S�m�Cԭ\���Xz�� By�fo o\bPb�P|�Y(@"`T��Xj$��o"P��q���kN�y�' O��M<[�U�����nN#���������}$`��]X#�P�]��xY$t�~⴦m��0=�`'G`s3�3EЦ�r q0���"t{DD�����m7�j_�����u ��}c�]+TT���z�qX������W�
�&Olukg�S��E	du��)B�K�)���]jh�١���D+��XQ"++ݞ�T��ɒ].�̜�
T6���>m߯abrÝ�;M�8���q�GȞ�^�z� �7����T]�j��w�M��
ʢcTm���e.@�Y�u�,�u��DO����)k	_��l��#�x��h��lǣ]�D��R����#�qu&��E�?�~�]6ui����S+�v����&���D��c�p�P'�.6eS�O�FV1�»������5�fu?o��o��R3��.��w���y�Tӭ�<
�6���}ޕ9��GS��b^ ��' V4�Z��)0bY ��`���8M�M|�RH� L�T���j�߇f'�=;�N0c��'ȑtuՋ��2���nE�ť��$�K�S�z�g�,U��	k	��]zt�^�"u��H�E�������o�օ�ot63��B���ǿ��p����XW;o�oR��K�X����uU=s\;MK�?��0oM��`���Rc�eP���XDsf<�/�S��vN�(MKV�@�U��bGe}��r��[{����a�Dn�ս�^!��7����/�~<N�̸��GLE��M��;��!n�Ē����N���'���y��7�چk�����8��_�������_�3M,��X@��Z���4�:�&�`�Sl�E�\�TБ��!�?b�x��.�hE+�z�2�?�n���V�h+����ӮTzw*�}d�nc���T�ܗy�R}x��Xy�ܩdSO���hq+�JD���u"�����pe�����&E���?l�^�ig��j�Aǈ .��x�N�D��C>j��%�h�stz����|��m���Y���0xI�KC�&��_�L��DET�֓O�V���h��g�
X����$�$�=���x�B뱯_�y���+P�JE�_��D�{���g�|㜘iҦ�SiR*f���NtX-:�6�ig�bM��9�8���	m Bw]�鈈&bcOQTP�'�)~��O�@e���E	[i��(7-�`q�*֝���Ʃ�'�v�{�->~6<�����.��9ʞ0�/������aZ�	�t���!I¥���먭�ٿ�N;�m�
=#F?����~!�۬ɚ{'iZ(�ԲEH���5��cs�·5Y.<�;~�l`V���e?	&چ7���Y�K���?B������[�5�$x�F���o�I�ŗ�����f�K�]/z [K6�z������%��L�l��5+�wU��e���<�]�(ϸ��D�ƾ��Z�j
������yh�¦>��C�4ѡ���m����^Ii�A�j"����FE��T��k�{� U[�/>�7��_���i !����,;���^� ^H�y^R"^��2M�ꋘ��l�Qg�J�=ҩ�.�O���)�Αti�CQK�X��d�o�O�~2?��е�JtS��0(�uɘ���r�
][��ov�Uֲ�gu ��we����T���z��G#1��������#,!ۍR�����UG���tߤ"hTx�ջ���,c��X�/��	�-;1l~bQȈI�즚[&��ө|*��u8{q4}�N�_���=�&�����#�"<�2V�#!Ө6�n�,��խ#��z�#sd4=�/K{5�As0x�����Pm(V�`��`X��5�Ujāk)���Râ��Ir	X�)Aٛ�a+"�{�*Tij���/�7)��XY=��@�,W��{q"��^��X��D肁SXXfG��xS��sn H�n�������ף�`&%X�����m3�EZX�?�T�h2��	ԾU:�u��{����v`��|�%B8���M���U}���X�9��GO���gq
�P�v	��X8�ڡ/e!A�H���G�
�[E�v�8R�5}�?�1���1CC:ɮ'z�~���SؖG% ̫q�In�~D۩�Sn���~6�>J��B����0A"pۗ�-�"����0s�X�b��*l���Tf3�j��Aɢ�t1���o$�Kom�lu��d+���(;��J}���bl43��
�&�%��og�;1ݵ-z�y�K�}I��5�Ɯ�m;�ȼ�8K9Y���$�"��4nln�)�U`��3��vBI����P׈����3_Z��: