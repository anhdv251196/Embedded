XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��߇|��q`֫�*���X�3����.���2�,d�Φe�`�!Z"���<碢w�D���1Ê{M+lt�pc��=0��s�x�
Hd\ysC�~/!�.˲����P�����7�~�t���n�6xM��x{�~��~�4"�3mt�;Y�J~�Z)�?�[N�F�o������m�d�����'M�+A`��(#���zW1w�(h�_C�-��ggPl��[&ִ��K��j�Af0���������nA��|�`����? "w����m�$]��ȯ�!���M{���Vnň���<�>$�����_�U�%"He��n@N}�+��/MRQ��Q�Q@m���y-G� �{�M�5�O�^Wu'�4��I�d�ۥ����'�2zDE�\Y0���)�218���m��.>�� C�T����#�c��U�l�Lv\��w딴+jZ����Uq`V�|)�&�6Dm^_�]������;��Y��C�*U5������TY*~Ob.�4�XE�tÞ��D�Na��+�}����(��f��iA��|'0`g�p��B��e��Dn�b���Vr���ѱ"}Q��"���� pS+է�̑q�ޑ����gH�ڨgv��ʹD�C��i��g���$��o�������ҁ`�˩;�gy�˜a���E��$y�U4�^���=O�����`�M4���!�e{�[d���D�#�f����wQ�Ӽ�u�,���<�H��`��h|�G��&Eyփ��XlxVHYEB    41c2     c40U`�_�R����`�S[��yFe��ĦW~O3��w&� /�Om`�5��
V���"��g�H\ae�,f�2�ůJm���O�5���� ��U�0��_��[�\5;���Q+M�>��B��<[�㊻����#�W�����U���^��������@�#�)��4w���.O7���7��q�%��V�s�m��U�_�?�np��@�r��[�+��֓E��� �7���Lu��_3w=��@7�i�NN�0����;F���bȑ��+��^�����4���uuv
�DI�g�U�$M��w&:gկK���ԛ*��+�J�u�Y��~:�
�]����s"MZ��Z�4h5	J=������En�	�	���9T�Q�(=u���n�+a���.˪29����7���{ټ�\g��^i�[)[�h��X#����䁓ZR��~�"a�ۜ���G�ѯF`D�Jj���rL$��잷I���_�t��%a�Ҽ��z\�C�)�Y��=�g���cEh�����&<��RPo�����s������?�2��n��}�X6V���O��l�����ů
�wk���ѳ��e�93^�2R�hm$w��<�'IȨg��@�X�D�)a;M�[�,}����<T��.z1 �{�r3sln��BNt%I�7P�0��aKf������Q�r랂��z6���G 3�]wA�d�2�h}F4�~�*�*ر��2��eI%5�uB<� �;"��C������o.��� 3-�o^Q��3��TUQ.I�f$��Iܣ���s��cw<�~�Lp�N��hl��RA��5`�I�3�~E,܎33���>ڕ�qq#>��h��/�]�X!�NB�øL@�l�A���ѳC�����40}@+������sU���Ȁ�v��u�Q"9�|JU|S�������I+� �as��x����bxJ�s������5�	��kSS)-,/�7I��H�Hry��5����	er9r3^�g0܋��ٚ�Ҩ�_�	���`]��H��#SNn��R����f���yt��������>?$D:������曳��ja���a��L���|�y�~����RT[��.��W�ҡh��������rCة��j�u��M�f���Ă��R�.��s7=,fK�iJ����븱0ބ싺ߌJw:�-C��g�hIdz.څ˚E��29�u���JKc��{]�W�^ �Ŷ

�Df~J���Ǘ,(��/���}��:q榴a&Dv���;���;fϸ�T�	S�3�����w�W��@a�������U�ڕOe������lp��p�#({=�g}�/V�v~�g��#� ;�G����]���K��  �R��od�&��4��EB��(Y��̨,�a��
��!�T+��k����%q����χ59�ӗB0G�(b��;�ґ����)yU���OM���\�a��͝�س� �S�1|�1>�i����k�KIو��#�,�{.�.�Ӗԑ�^*�P�����Bm� u�W(���f��V'�k|����m#\k�Om�����;�����?��y{wD� Yzes�V�߂�m��&L#""������2u���GɴG o1���G`�W^��ebe(dTp>���� i�?w�d�����Cܙ�{#l҉vo$���O,�y%�٠��4��w��B�m̱���ZG���C���h��-k��v]�[GF�|1�i���@3��QL ����zSsw�<��`��3%K�я��O���g��\_И	���Ι�r��A��U�z ��{��2��\����֚��F�z��>$!E�,���lAVyM���u��Lϕ��s�88��Qd��� l;��Ҩ\e�5����Ma���$aȢ?��K���|I��y����_}�G��cpѥ-,|�@��봛_��ۂQ�ˡ���}+�ɰ�{xR*�]I/ގ�[�~ܳq*�M���Z���S�E{�IVpo��6�u4O���t[^>���M
GO1��`T
HG�dyFć�/2{�� YTZb6}��w���C��z��lB�ܿ�Gw���mz-��mߤl�����}�FLe)2gr�cd2�s�[~X}7Lv����N7\��(�N:d��1U!)����a ��gf��&�V�M6V��n_���6͔��e�	�P/E�4�z�D�߈!�����H
�=e�X�W�h���K�����"�Vq�����"���?�h��-��=���NO9�L�B,$y #��0�����(�d6W<�L���m������䤹��XjI�]�p���;�R+�s�~X� ,��pV+B�#&�ׄ�|/#u-��|i�7VG@�5m��{U!�s��3u@^D�{��dHX�*�-��o|^K��{p�=H׌�[�r�\2G�q�j#�V��������7?�����?�\4b ���i�$�NQ���̕b&r4�A�[�D��O̥��e�\k}E��T����^�P�{�~*�y�L���"���hǺ��rc�j�d�:tT�g������#����¦�}�8#r���,�6R��SaW�I����3V۷#�8�?g%�tcjaqݫ�e5Ty�L%�i@7L�L��Z���}�t6��b���-��6@{o�OK��Q�΅`���&,]��THJ.��.~M&8�Ց��Dvb���_���6�����s�%U҃��1	3�+�%"?⵫ܤo��G�pxu���/��#B�a�U\$�*6�65s`�5����^Ύ]�c�x<�!1���6-���%���t������g�N�xj�%�2�k�|�bX�6���V�gP����i<�].���(Mo�q��]��~" ���Ht��6h�b$�OQn@]�X�o���9�����]e�� D��;��t�2�5=[�Y�sY���@�Kߧ�Μ��B��f�n�6�<��~M=:�a+6r]��ee7V=�[�($�42�MT{X���ꦰi��XR����H��䗵̢Pq5gSX�Q5�=���p}d����6�X'�S��5���� ��v�>ߍ�e��\a�7�]���r���ɒ{��w�X̙/^�/�F�JQ$c3�w����������HĨ%o�