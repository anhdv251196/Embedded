XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����K� ��9�@> ���A�U>*Ʋ.J�n,� �����^�v�̎�6m�Ba�;���E˅�z$��kE�w��]s9�s�Ge~������L���o���mMc�7XgS-k/�!��'��q��m�
ɴFꉻ�����n yy�S��Q���o��K:6�\��мqRph���bw��$��*CNMh�l	ԗ��P���ᑳVv�0o�Ĉ 7����e���ԣ3�=u�^��Լ�`4����"�>}h/ݜ)�f5��<3�˔�C�7yw(��Ǟ`�(;M\��5jʑ�Z��϶S���~Т~�qpϯA�� ��N;_p���&+<:�l8��/����CY�E���Lt�`�-Tu�H�A�P:+���;��@�-�������5OCjB)�����Oh�TOG�5�~�����E�w�e�#`��䔺o YH���U�����c"�
4gyO��=ܹ<����%䅪,�"ڦ�'Ih��1�����u���a��i=w�os0,�iR'd����RE6��"sw���b�����V�)�j�;���l���B"��؂
�|���	���_���e�v�����*H���M�$Z�ƻ�"�K�����5c����|!�����2����Q���?y������y�d�U��
��|yt�A"�Ƈy7j�6YK������.q�
A�1��SeM߬������>&�6+ik�9ɞ��b��%�&
�Brڧ���P�a���͂�4�5�̶:o$bJ��XlxVHYEB    1cf5     790P�-�{[�QL���W:��1��'[�z�����O��xxf�
�A���鰔oL��^�H�-J�6���%fn�HN\	��r�p�,̋�%LG4�@�05E��%��3����ȽJ�c������>��F�+
�$u����o�L`MpD~+���� �<�ї����2�0���l��o��7���(8��r)q���,�M`���e�D!É�S��Ҟ�H��<�@=#\�����1b��1�b�o�`�S�HԳ��ä�V	N�"�j%fpx�����*l_�wH��ZT.���!"��)_ 9�������C/e �\{��ێ<�u�v��0�{�O��Y�h�{b' ��f��E���;B�yšUT�]�\V:2��D{��5\N��N�%b��u��6ݤ���:l /J���6g�����:;*�"�L�+]$"Z���3q�2���/h�^�Ȧ4o�=��'�WZ��ŨJ��;H�=IP�N8�?M=b��rK��v/	*�{����:?c���O	"����'x���`����c敤��&6��vԲ��"�%��6@��7gpW���S�ӎ;�6:G�������s���c�dҁI%]S��%�Z�P�ri�Ƥ�{˒0��(>�����1�\ȳ�G���SS�U�����'�	3�\�i��GA�B��Oňq/V&F�Z�c��b��c�Q#�;l'��> `�6�-�,���l���mn�|W2g��,�Q?���V��J�$;$�P���7�E���^K5�k)�wX�0�Hg�C�7}ĻO@ˏ�э��a�d��>&Ē�ǩ��~m�Z�W>`@��2f�e��{��7y���_
׷��5-���E�u�`1;#v���yI�}쑹N@P�i��
�ln&o��sw/ݡv�W�ֳ���`bEB�G]Ü�]�ߗi7^���e����<L��Ez7�yOj���wF9���_�G	/�C�ho:�����.���/>����wf6d;e�k�:,i��z td|0�b���`V ��6����2����BV�{:�n��	ꔌ37M��蠅�KY8��C�����T΂��3/v�"'%���P��;�t���l^	�����(|g���N��+4,z�?+Kx���4���	�$5�~���+��_}�G�pOJa�&�p�2tה�(z\r�!9�c�����	�:GrQ��t�������S|óӞ���֡�A(�֓�K�W������J��y[Ni{�^�'�/��	�^띅綴��jKm�l�k���N&�>������e�Dd����2㏑X�Y|
VO�Us0�f:M7�%��Oy��wfEZ�gt'���K�g�^d��-@�y �}�L
=��G�>��vd)��(u�?v�.{��5	pX�&{� QMܧ��d�"���)6�O�qC|���}�.�#V�Q@���8�L����T�>��A���y�Q֑��8�iu�|L7NA�?�[���f�/��J�����7���	i������x4�������o�a�[w�[��������5���{��T�Z��?�����}�wRM,����	(c��b>]�h�X���6����N/#hY�a����u��xزH�{�p��K9��F#��j����Q��:�k�x��^V�0=X����KP��JOp�_d;�kn��v(�v"����֖9A?�@y��V�z���zP�U)���_��]E��`����Xg})=܍m���L��qʝ�u	2l��<�̯�,�e	��֢5��J�R�k�%pN�g+Q��(�3��s���p:��y61!}�S��	�k��|�(�:�(�4�X?Q���є��Xe{��#��gY,�B���Y���3"��Xݫ�&����.c��1鷍�)&����