XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��[��w7#Q瞄����?�@�j\8�r��_�B���e]�DK�i ������Y�g% P\<EZ>n�{��&P�s���sHX+[�p��SF���������P�������w>/$�E�`��Hq�VM��I��J.:���گi�������W�0���M� ��{hɊA�&9���s�g�l�yU��ͼBa�����Sq
 j?��O߈��l�6�Skg�D�3=��t�+H��jT�_��d���n+~�̺8��J2��F�5�5vk�P�S=�H�1�8��.j��f0ن%�2��!�!�ss�c�RԂ�Xu�#|�eWKr��İ�u~�k�ʔ�=�Ig�h�A�N�� � �etb�,V������cέ��m�E�=Sʚ<[�L&1�pR��Ć�U�6�A�0�#̨K��#����6#Y�
,N��=K�I-��W|/9Ω�	��\�kP���J�E}AO=J8AkمN$�'%������^����0&�?1Va<U�`ш��/�f�(SPfދ��5:���7�#�PTɜ\��f�I�)ك��ݡ��E��tr���R+U�u[H�U��ަ���?юM�(A�nl���w,�%(�%���m���q&�>��J���c@Q�٣��4r�����.�E�����t���" ����{��}�9�g'���S��Q�U��I;i�y���Y�����=�|u-�wW�6���*V��#���/�I%<��[r���щboW�ݹXlxVHYEB    6faf     c30g��:�����!-��C]�],�s�vd��;>�/[��/����������'�*�"HP��b*��C]��������xq����#�/�3J�f����I�$,��iy��/����,�~�
n�)�{�n�?��[�>`(��$7�\��Ȃ��t�mr W�P�M���i,4,�7�W���"�����	*Vf"�D�J!���Ԣ�,~�O��Un�u�T�0��L�-E-���ފvqF,%��������E���wmRah�C7e�@^ޗK�pR���j��v�(}x�+�9@U %H����>��1� ��V��=��I�7BN辘�njZM�������#od��v�EE�׮�������"�:�W�,�k�t�r�t��S��W�xbd%u��h�Y� �y�p&�,��B���}�����`�����c#�/l�Q�Y�r���猙/�XYm %����-�`������@�DD@ZI�M�2�7�7��jg+�.�T����K\D@��r�G��^��:EJiJ޵�y͙{�<�)�繻�ӽ,���h�8Ǫ�/�Q`�U��"���K�|�V�q����k���q�m�I��r��c�rS��^#���Ё�[;�f��b0�W{�YC�X7&	�FY��sgY	�.9��	u�dG"�k���l�~��(�������Ay��u�z��*�@R-��%�*��i�.�0���!��~\ls
���N�Eߕ�k3i�����Z�e=h����k�rTݰ8�1_�|vO�����;
\b��X�Q�X&~U��\}�6K#�ՓA�%^u�T2-O���[}��
���$	���ޅ0��b�R���T�%�X���%�VXW�oT0���g)�κ��������A�ƃM�h�Ư�a�C>wyЫn0!j��+M�rum@�v���a��n�]��'s��D�d�(�N]���96D�#G��F�Ĭ���R�/L�OF������T.��DV��&��W�٢��,<I��5v�v��
������]��K��!����Iњ2C�^.e(G����uf�@�^���a�h�F��m��}����X�H�RN�n��uB�T/H��~'�/yPAT���̎��[��GK���i�q2s<�~�}!�����prjq}�95���}���Y{@MO�J-��n�X��7(�4/�\��5��Xp�8\e�[(�F\�A:�7�f��U�֑���U�d�7�/r����D��Y??��̋�ss�h�r�&^�S�%�_�+�J�Nu��~�e���}�L�<��u`O���:�G�R��lN'�J��ڳ8J)Hΐ"�Rv�垖t������D<��Mh���?9Q�H<>,&��^��	X������6�|�6/QQ�i���m�ku�^	{�˷d%7�Ԃ1�vB�`���Ρ�D�\-`e�@HC�(��)\WC�433����{v��ʢ���6���O���3��8���6&8%�YΛ���S|�i2J��kna���i�b���H��h�<�|�7����Y�ZF;�K^�A�����]vXؾΑ�.W��@\p��lJoRSx�'	�\�Gʷn�4sI�EM�)���&3����g;y�7i�샞F�Zz$bs��*���Bh�)������B��	�?�,ӯ,���)��o�s���j�z7C����Bh ��
7�[��I~��E�P3��./八tw��dյ��ӡ`�=Uz����O�__�X�>��j.�w�Wk)��u�N��0%���P����y�e������If�unW�|tlN�àGrp�ݘ�RfI�*&�,X���*�@���j���·�4�jo�C��Xض�M:�]Վ��ݥ�Lo��[+>��v��+U�h��=�s ��@�����2�E�`��A����L�3D�laLФ� ��1�ݻ�}��[�6υ���[vًHe��(5/�B^�����Z��;	���7��l�����4��*�!�ҝ7,S,Jr����44�D��`��;,��%�8�i�z��A�]Kh���N��>�fD����m�KIU/�rq�EBAM�(#�2��{c���r�t�1!�7�]��Lς�,E$W�u��疮O�O������ n=�8{��ۇ���x���6��3�5`#��AO��_[fhfAgK��P�0�<2�{a�^�&}��;����5
{��%�%V��<�������I3��Z�G�h
�\�-:`��RQ����^Fm�d�c_��8p	�<(��s^r�I�}��{���B�M��/]<�Q��y���l_T{ԉRc�]��U"�b��Pw �P4��������‣�Tj^�lh8�| �ʒ(V'��1��?χ"����3����q�M7Ⱦ+�H��\����4��it� Ⱥ�B�b��1x&ѝT�e�N�����x�'<����ѻ���_�c6Xeo�������)d�0��7������]�!���HMt�YW�� e��р���g�����ۆ77i�_��6�����ע�^�EhN��i��&�zLU5����2�l헌��t�{٩V��m\ڰx�W��b��� J��7���v��f�S�R�,z�y=�����ݚ�����U��I�^�a��	�s�������m�	��c4�ޜ
�6���fS����]��������w
#���9�D:�$�9c��~F�L��qȚ��`�Q���eC' =��5����!�q��R����~���I5�{Eڡ��`z��xہM���#,l�3s���a5	���kYr� }�G��u8�ML/��4�8���"�D+�E�E�����+�������珳��9�X��<L8:�;h����d���>`�Og�;��VI�=uo����)eC�F����1v����Jn�(^"��D\;&�����t�|~t>E�������S��[�0�)9�ޒTWl��O�c�t%�bi�
`Q��T�e~jf1��3�B�F�����jH�RB���Fj��O�����ZS��1eM�'v	�5��� ?�.^PJ1�i�@��t�2��$<�*[u1HZ�_7�tl�\������