XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��#�^i��Z�"�-Jb\�5�~�]<����^H�/|��if��Hn�̻�K��)���0�Q"�m���$���#�,���&x���x�7�-;Zt>� ?Ws\��o�i�VH��.��ȔPwaXzWgA�ݪ�3bפ�$��{�/7����6ƺe	�E����i��<C@c2y9i�glm�U�kCߑ�ʒrY*�O���D�1�Ԯ<�)�CJ�bVt�%t�@:{S3*L
�>�!����*��߼�k걿I5o�?���2���>���S�W��1�JC���n�|Y>�?jgBӼXX�x�Up�o�G�*N�Ǚ֭;�ș��a_hv����N�m��ʶɊ3�mhv��?�#�c�����	�ߊ2zӧ�����c�,T�+W��xp���?<��1�/᫜?�X�2�QJ>H#�ח5�G1"Љ��ۦ}?e��ŏk|����/���1pYd1=��U�]ʠ���Â�z�~Rn�g�й��rI7z}e�������Mܘ��aC�q�7vV4���/U���G^�j"���@r�vΕ��4u�so��6'����+^D?�N��2�$�B��h�ҡ����������T�'����>�����1����z?��]��,���}v\n0t��w���q@ 'yv�ۆ\�E!�HY����if��c��Y����6���=�c���1�C�QL�/�2s�xk&gm����5ۅ+B' �Q�O�M�p��j_��������{bMXlxVHYEB     b05     370@d����Z�?Lp�U)$� �*J�ۙ���q?m�-'�
#Q�I
��6����W�ܳ�	�"iI��(���7��V������+������m�
�6uE�#��4J}~q��y���JQyQ5��(3���fz6}�� ]��[�m�u磰,���pԴw}?*H/>�C��{�ٮb�I�ˀ?������}:!��Dw�/m3��
N�X���Z������D.r�¶�Ƒ{;-R����*�X�A�&�L�\���G�`�)ɷ�N)�pd��&�M���F���^X�W�-��Aɧ���C���q3�GJ��IS P�VNT�j�u��)>otY��#�m�إ��Q�-)-x�/K�����$�ތ�W���:��	d��TUj@���"BO3�ަ��@�O7xǎ�DP��1Sd���=�$٣n9�U\���|�5�^�8��=�^-f�L��������O��׬x��Y/�yQ��hP��YOaο�=�H
@K �X�� �Cѕ<���ڒ�X��C��ڜ�}��bCNZ�i"oW�w�=[x���9�l���7�q�x��U% ��k�ξt������I��Z�z��^'�Z^�iM3Yӳ���`�l��$P�	���)qn>�����&��ے�krȾH�T;��K�ͩ�+apy}d�'YY����z����OH��U�;�����y=g�پ� P6�5��E�9��!}��V�b��z� �3�������1�pM]-4&
�\?d\�A9��g�����NA��J�%<,�'D B'M�~YG�����ϯ�=���1�눁h�C���kt3�Os�Dy�u�]��`�©�O��?p�;�#�_%%�;�^����9�