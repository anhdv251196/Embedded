XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����??�p�Cb�#���I�#^Y�Pw�Z�\t
��{�9�(!�#F����\�5cw��"�;� ��0��'t��������j��Q1�A���y��/�R�~�vf*�6ܦZɅ!�%+K�q�S�� �W��>���@��`޻�=�~�x�z{4�Z-���ݟ�d��a����Vt�]�P;S���d�{�ZG��La �Ah��"t9o�0�X���-_,���h��P׌#�=o�4����н��sU�:/U?�癥 ��
���e���C�Nzx����96�y��p����k�£�T���S*�#�
��R��;����섦u	�����b��PgURUN��mB�D8�D��~����5�e�%6:�uo]e����鱃�#(��c�V��L���L	���	+0 $��L���)p��b�/'l����VR�E[�6w?I�ln�neӳ:��T���l��|���*o������6�ଘ�u�	��r�,�oEq�Vޓ���g��sD �%� ��Y�anm��Yʲە�\��b+�lJ&�-���`��#�#�c�1����PU

��?G~�5�ɵ4���6<+�k;;���+�s�s���c��zߞ�(�1VP��y�UUl��Ÿ0h��� O�S�v��'�#�)/��-�ᅥ� XH�Y�g,|{��.{\��c	��:y
��mM[�&��D3r�NR�!��O\/�Q% O�}�W��Gz9v8,ɫ�tD��x�
��Cl�?@XlxVHYEB    156c     590�䌡q9g��W�N5` Ӡ����:�NU�$`��=ʑ��Z�~���:�+�p�O��?Fa��Ḃ�'��g�6�j�K��W�4��H�x�qF�c���,´q�j�����إq��7(����+����T9�h����s�+�˱��{��t��W4�ﶧ��h�t��t�7�L��SET|�`�\'z��>��ֱo��8�k��K�҃�/��݉O�5����|UAe�Y^FJڊv,L�ke���m�#�M�0�������D7��B���N���UG���ThoY-����_I����@�Z���((^��N�b��wO�Da�����Ğ:�K�6�!�|d�I:~(�mϸ8`
�����Q�L��|,%�#�<�M��I.�Hk���إ�A1�|D��4�+�Ed&U�x��Ǿ<����9Tcś*f:*npN�(��B����T��]#�������!`�]=e�͊ =-�Y�̆�~�Fɭ�v��UҀ�v�b|�1h��>�4ވ_�,���,x�̰Z:M�e`R�缒ͫ��Xkx묉X"�k�Q�ai4�b�^@d9]��G��H�g�@��E�f���tf"*H���ꥥP�^p��k19F�
������;�\�+���7����&	�3��&m�\g�mGŻ�5v�2Y
�"�&� ���Z�ĕ����7Y�ӌJܪ��A�U�-�x�g+Pi���"�?FW�Wfү����������'��C��0��ɘ"�又7��Q���hh\!_A�H�}�j�����SAL!�f�ΪJ9�W�z�[���cJ+3#د4���f�w��
T
�����d�����PƣV �Ԯ�K����{����	w�E�\��u��T�4�ma�X\�h��l~:T�z0��sw���7��|2{�ʠX9ۼ������_5�'�2�w�zBy�ek�FE����,T��:�L�ѭ��c�u�n� ��9��W�NV��A�&���cQ���f��/q��	�	#.^Q�^�4�/����啈��&��4&�A��������A��4���;K)�3���;�n$jID��c�?��c<�s�Mm;6���� �/��n����C��6f	_��.�8r�z���L۔�dc<S�s�D/���Z�K���/���
-�}�������ǭ�ș�(��yyAl��� 9���*h�9���'�Dy���o�?��î�X^�BO@\�O5WO�o��a�7m=H�k%G8��s�i73��e���j7X����(uUqHmz�"�&̠a��G���6P��3P���8�oh	d���[$F���Gr3���E��$��Za�Y?DJ.me%�L���T�0����ٸ�� ���M���+ex������,���4��P�Հ��}Y�(<#cw�M��/
��