XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���s=���WY$+w��В�&ˈ���l�.���Y㏙��Ŧez�6�-1��Q���i2�	4����kR�g�w�(qD/��+���)���~���v͑W��<��<���͞a��,�A�q_6W��pg]��v)�	�������	�"Sl�h�1�<:+��T�ְ��Y�82=������$\q�@���������kjؓOV'����H�"S���H'_b��^��So"�v$��c׌	��CR>�:8H�J���I�ң�.V��'�Z�������F[�V�=5��0Yd8�vz�6��:a�
���E�/BE�Z�<�a|��o3Z�c�	)��Q�8�m[;�p1���kRf�KX�ڋ�S�4�H$1%�����L��k8�ֿ��G��_���D�n��g+���_��Q�A?B�!5f܈����M$�oJ/E$��0����Zf���:���OP�^�����^�>$�'�����m��y���Px @e�"�$��%�O� D	�!��_|a�@Wt���!�P|UB�y`�k5�>i��mm��~�wTYx�|�������?�����7����B�<+��VD5���!�W��,!$������'�~I��X-�:8DJu��Ǥ�m/sX�X��/k�>��<�ZX�����R�/Kl�: ki��*����~.�Q��?C��SQ�q��*�:)RT\�9G(����Lv�^��Y$���$�B�C��'&6���-��1t���)��x��O��XlxVHYEB    5a4a     590)2�^�#"��fD�������C�[�6&
�����"@��P��`��G������인�a<�q!"�:7|�N��8Gd̢J��O���|)���ÂH�]�\�+��6k�kG1��c}��|����H�t��O�E��ݝ́���a����{ek�b2Y��(w��,��2���X���h�(��GB �_}��s
N��0v��n/����';�����p�5����`���e�'������A��qe��+��!�w3(�Yn�)j�s��b}�#�7����!1>��L�F:���0�����B����xZ�?K$+�؟�~�3�X~ܠ`?�E�Q'*���%9�3�Ng�MW8۰%�&�ٲ�l���q��e�{���J03�? H�N�2���X�Ur=Rc'���aю�������7.MiwƬ��"c���##���e��hlk����! h�E)���,^�?v>g�D�f3����0O�����B�����ʲ�<[m�G2��u��2#h�J�.+�G��ޱ���zP��ɤ�4Ggz����kGL�9�W@�1��Do���lƺ9��N�
�=�Z`e��1�ʣ/Ą�q�i��m����(SX����ߵ�_W����QWG��T�A@�L�'kS����2���h��o��,zz�\������	�L��~����aL��"�nfħ���N����eq$ȯ����Nm��&�'��0�6F�Or,r�6S�����11�O8��� ��˴�6�2����smw��3���P�m�%��C��n�*O���3����_���'Y��$��{ �}���*���_8�Q���ײ��S��Es-����s�	���]�;@H!�n�(3��H�*��	~l|�9[n�����Qwu7�S�	��)������m�����5̇��I��<W>�&
���ϵ��'��.�@��O�%[4HW7�2�*A�V�{p��Ǖw�L|���_�|���d^���en'>�h��ۨ��ғ�� 쎛�����9V�.`�Ɏ�����V	�h��Q,K�%
����TJ�?jv��
���x��ڥP��j��ȹ��D��m��e3?�t{-���~�#�<�@���[jĠ�v��1=��LQ,�(�pP�ʇ�h��WR�u�Ѝ����R��X�VO̽T�,���$��`�Ǐp��J�"�BӱD;D�q� Ѕ���tz//��P��f\E��l�_�Էy��b��~����3����N�| �|M��Z�B�jgЖ�6�@���1<>ߑ���+�h-c �x�=y]�&2���a���N�4{�K'�;�����=kg�X"�5e� <�n�`����w�#9��DL����>���R�z|�(�幀�Ɵ3��ǩ˶��w��-x�p�&]�0