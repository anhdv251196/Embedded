XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Ђ�<�=vJ���V����ҋ� a!N��jG����%{ N%��V�უ�'Z�RqE�g�T�=ƅz"e���V�./Hn��눹��	P�4G�5IDVΛ�ɼ�Hb�F<�1�+��v�s��q�yZ�^4g]B�S����t�:O�̫���� �=��icC�Oh1�ʟEOqb��{3gm���\(�jn��QO�T���n���R��1�T��hj����B�UL�S�D�l:����5�^R|VUh��tЂ��m��4b _��Q�3l���J����Ix��+��a'��$�B��Z�$�=K��ʹ��I�jf>�|�����M@c�����{���%�CWTd��a�?^��l��@TZ�
�X>ߙ�n���kr���M�(�1�@��"��V ��ݡ>�h��+��%j�A(�"`���ZlX`��*��8�}'Dh�AN�"�@����ػ�V�{H<fw���SK����A �qu\�PP���[����Вf�i,{�g�pI*��������+p��#&ɸ8NB)We��"�{>���zH���<��e�^hJ�绾J(�����r�C��'���.K(�pZ��bU1祈�������WH��t����c����Q�/��8)桎 {G�|��q}=�?��$E��r"��,������@eֽ�f�_���2i�;�HH��u��i@%�ݴ&���В|�w�`%���Vj3ϕ��_B�/���o�/fm㫄�D<?�?� Qn����DXlxVHYEB     b35     3d0>�W֖ӥ8���l�^ �w'%a
�)�ҭ0Tj���Ť3c���&���Lzx[��1J���i{�T�q�64'�ۤQ9�{'M5�(!�Y�７}gf�ؒo{��u�2�}ը3��W|�zz"�k�� De���;�Z8p�h�<��д�?!Y�-4B�W�8;��DI�M��x%d�߆��d��4&��R{��B|�b5����_CGn�D��>��b���g�0Nmj�7�āO��0�<�6W���П�^��T��qp�ޛ9�7�~(<g��hC2�P�p���s
j��P\�-�W���N��y��J�tXXM��OXC$�E2��}�|Dz0�������9:Rpg�[�s>,�!�聊��cI�;�i$#��ji"%�x����,�x�qʢWjW�z���$4�M�?�jC�0�v�$�i��^�!T���V.5X]ϋZ��j���	�%`�޿{_y��`?�inp�ur�taz:�C��Z�lEAzu��"�+�	�O��V�^��u���K�r�[*B�n���dPA�-�yu��{��lj�uL�ȇ��(#{������=Sˮ��d���]E��s��
?�g9���mwQ�(�%:�h��XB�)�HCb��=�!µ/ 3���/�y��g5�<�|$��P�x�!K+�"[qo�Z��܂�����U�Ĭˏ�;Մ�)�5۪rȷ�z0���7c%Q���ۣ���7� K/a�t�)�{A��Sò%ay\���0p�j���m�[LWڮ���3�b̮ݧ$���9,���ο=M6ALi���=% ˎѭ� �K&_��g�)�g �]�Vg=ȸ2?�P-�9�X�L~�
�_��j�k c<�S�����݊�����?�0��� ��־�C<T9 ܴ8Öp�7���}��߇����c��ftz{�<]��
����>F�|���<6���.-hy�T���k��J���c�