XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��gc;��7�U!/j��J�Y#��U��oi�7�����v!椂�5���:�07j)�[,0u��%��pj�#��ԝx��n��b�G�/iw���?�>�J� m:���~aM�B��u�l�{�U�u���]�ESr�㉵�l�?[ld��x,T;�V�-�yi�f訚V�"��^�+z�67υ;��b׊ d/�>f����_?ߛ�k��"*P펚($�t{`��i���C�Q�64��	"� �`x���{v�]�:�9�E �k^�;#$��7
�v����/��+^5�F�d�1=$� �5��� �}��մ��෍�t�q��8�uKTʸ�!��(j�<d�Q�d�`�h�Q������zH�a$Rl]����
e�x�T�܍�n�e����_F#�G�^
p�5X՛ѿ�[��H�s@zn ���Yn��Ԡ2��iE*�����W6����Z�;ӱwZ�i.[�W�o�49	ek� � �ڣ�T����<����_�&,	Wt�<���	�&��uf�.�����hea�F ܗϹ �N<`�́.̺-Vt��ğ�݃7)g����ě>��n#�֏�i�>���O��i�sena�^�O�����7m+Կ8�����4K�xȇ��o�z�qɦ'+���r}K>�7�J�ހ���+<#@��"lJz�6R#!��+��n��$����5�By�3U��K57[��+��دA�|�Rc�v�1_k=]�"�DCZXlxVHYEB    1d53     7b0b��$4$1mGҟ�rG�̨��/�XMVbT��(S��Տ9�Vą<^��߆��#m�O��	�(�tCG4	F<>)�3���ϊ����Q����2`6yw\���/+���B2m�(�k�.������q�9�D����MJa��� $md�_U�^�M����Y'���"����(:�r�_���Z@8���oF�MĲ��N��̵�������bq�,���"�m&2�4�3�	�%���_���$����)Q��뙨����"�k��ܼ�͉����5����F�CC��z(�u��hN�T�<`|_Un /� ]�<���?E)4�,hh#y1 
l�-���z_y�+�%6�3���xu 0���vq���)�Ɠr@��D��ii`
Ƿ��v\�N�f����`����	��W]�w#ȡdZ�ߴO�@\/�"�b��k��3b1mĦ��ᛸQ���~�2;<�zٝz��a����Wv!Ŕ�Ո�W�����Ĥ��j�\,�����ʑV4�%�P�D���(��-��`<!����Z�I��sK��ZG����J-08X=�|�Z��F�v����r�9�a�mu~������k>w�Ei����x���1�BE���η> N�����C�z5����W�'>J�7r�eGA�eG�֩�=�>{���x�}�쮼�y/�7h_-yJ���P]]Š����Ns��Z;��
��!�I��]>%���%c�X��xS�&�cs�Cle���Z�0T�.h�"��aU�⣫%�Z�z3N�b� ��~Kk���ɃdѲ
��b����&>��ڈ�*#���[(Q��r�U�rY;*��ɗE��� .����x�fNQ=�( �:yA��a�L����yD{�t^5>p��K��3Nz�m��g�N���c"���b�?�!n�ց.�d|֬� �PM����`�'�I��]�4�WLS�����6��?)�94���f��yL�r�+�Y�Y�*���.O�)X�4z:ԝ��I�~�>�t�|���]�,PO0�m�/�n��b�
!qv�#�狝�sz��6B����D�YW�:p 1���$.��b/�QQ�����[�	6�h(���*`e��m��]\B�^�z�-]�������sĈ�=�(�&�KG��6�d��6��Df�&{�����ϻF�Jg���ɇ.[��/|	u�L�.��2��R!@���;�NE@?Hp��"��o��A�a>	<�^�W~Z�qi�#� �e_��]c�z�����e�7=KŞ�e�@U��qb��O���f���ߒͼ�?cR�Z�u=t����axmH�vD�w]}AMCmRV������s�MTrpZVO�T7.���b���ᾁ�,�I��*�
�WVӋ�p�/y9M�gІ��� D��3�WI���o}�zae�g���/6��xk�im�C�h����^_�^�	����vs�;�ޚͬ����_������	�����|%�|��۴�?m��&N���+y^������>8��0��;D�g����|y����+��'�
�i�$�����:�Ѥܳו�|���tx����βx�� .w׸�aT�Xv˟�m��ϸ�aꈥi�;���>qx$EWi��b����C�'p.x8�`��jZ���"���f�a�K�^}V��r�ۑN��p�|m�7�
½γ�U�{��Y�Wl9�$U�	Ao�|��[�r�򓣆��	��}ݏ쭕�X� ��:��G]ͣ��Odeԝ5?jl�5�y�De��RYja��������|�����3�)^�.�-�B���Z��u��u41��F4"��.8E)C�Y�BCu�^T7�{�7Q��(z��醿r�+R/�.6�񇣮0p�����1��	2�n�.c����� 9�Q��R���L�LX�1'�X��v�.^�E�T��W