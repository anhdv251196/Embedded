XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���T�t��d�\s�E`߅��)�����X�X�n� �[�ς�6fm�湀��d��	i�5��aZ�^O�)K���vB�羆�jÙ��v<hKO��~}��¦Ĺ�e+���%K-��ǰ�����ș�$�ڜ��J���h��e��o�$�k+�(��Po��x�f���O�tr����cG+e��A�c�����R���Jg�K�_oyEQ������@s�W��kw�N6'و�����e�ey�&("����mN�G�'�7����s��$~��n��
�u�+*&��"-J����<���hm��E�|s���b}�sCN���P�ɪ�t���?������}���~R�
�RÇ\q���*kb�v|�<'9�?^�X����]U��)��h����3�fػ�M��c�Kbo@���� 6������e�^�� I`4���T|���轐�Տy�o���Ip-8 ��׳�� n��%[�y�����@@]��ކ��Q����:H[=Ξ2hH��]ٕ�[�Q��7_��N,P�J4�	c&��@����Gd7*���4��}�
�;Ì���U�9RF%����O	EMX���:�o�R��4E ��Uh��)$�C�����\X��	&�u��g�oW�Ӛ��i.�_{�P3�qrT�Z��?K ֺ���b���~�겨���xoq�)�IfH"fka��F����R�_<�刿�y)u�T8(c�vF���qzE��Y�5Y��~~>�8<��!_7�ά�v��XlxVHYEB    165c     400&�p�6�G��[�Vx�:zպ��X��sR�݊>+�q?�Ϡ$ c �j��8�[�r�\ ��؝td����E[P:�:9.U�� 5-�f�T�&qsBr�u��LH�m3t=�h1�^G���m������2�
"?�|(��A,rD6nT-č !��(�`���"�:����/hQ��;^7=��֍�5雎����kc'V�}��U��ދ[e�P��̞��;�Bl�.�W�����VG�x�w@#/S�M��y���I#�Ӊ��A��4N��a����3�~7g@_��w~����r���[� :�)��}�FF�]B�$�w�#Ӣ��)e���I����N�7ez��j�ԅ�[��n���V�)���K��
�9�^
�VC������vX]	�<��ِD���1c\��,���Tq�C��{6+ݳ���5���s�U�Ŵw�-R�AƑ�e��	��9R��ϭ�v��z�T�� 0Z���I�K���@��f}Ź�m"��1����ظ73|(�������Vq>��~��>�E&�^"��P.�n�آ,�ܙ������5$�m:P�������A�s��/;�e�3�n��,M�a�T�
���k�1�$N��	2:��#�@��I�Z���0m����6!��B`O!�����r�R
�KSP��e�nl��Np���2X��Dͨ0X]���;N�f�E��� �xv�Dɭ�P��#^X��n���L�kH
�=��Ů�D�?�Z�r�咋|��B������D�4�]C��n��Yn��:���s/�g�X��N#���0o��js�` �]�O�'4�$�*�-R����-<%�\9{ ���}�KO$ӝ�.7)i��~d�֫,��I���A���
3z�JuT,q������4ڧ���DRT	�]��Њ|g���H��ˏ�B�D��ajt���!��>50Bz��==�=��!�:�T�%,�xT���$'�mB�"���[��҅�\cKރu�p**��