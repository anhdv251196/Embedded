XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��b�b��B���d��j`?s,m���S%T��i�����x�R����t�dQ�ӁK��f�"o9����t����əa~Nw��ʻ��:� �/��c2�@�=�o��]��h��zL_�f��ᣞ7��46��V�ބf/�Pܤ��	��N	�wy,�
��D�}[���XK�U\>}��y�h��~Ͽ-�$>���#�~��dw�|/�C#[$zL錯�W@;��8���cM��;,�g����U�a��^��8h?+��
���6s�t�O���Dc�=��j?8,@��ϙMT���4v&��]b�V�'9��Y�u�K�mۚ�KzĚ��qj&m�d����\hf��ȵ�b�C������	��0G�/�x�d먇�e/�V2if>�{��$F���;��Y� g?�&蘊�k��^�G!��9�_�,!A�1'P�����cm<�5L�<��azR�8y�N2_�0����]a��K
 �e�2qf�(!��L<w� A�P�wȼ"�)��+�wX�L�ѬTK�8�p'��t��ݴ�O���5y-��O�]�d�B
-J�%QV�;�j�7��0P�g���Fh$"!���^�Y,�3�sU�����˕՚%��(X��.̾"!�>��r�6�Oς]th�B��=�k�搤EB���wr���ȱ�o	��ʐ�Һ:#�+��hR��o�����a������M�Y7�BѬ���߀�EK�R�?ao�����!���M������1�d��XlxVHYEB    1d4f     7b0��j���IlϘ;Ѭ<�<y
K���~�08�SW0�����H���-kH�'���R�~ަ�� �A���'�`���hE� �|H�t4�C��8����h�{Y2��
Ј��)�~��T=-z�]fޤ�D��8 Q��U��IM��g��+=�.~�e��5:.��v6���Yά$=�*f�ָ���� ���[9�v��h)z�ܷ�D�4���&X���v5oGĔ�Jk;���a��<��rɪ�h��G��Ϯ[�L��5�[�|�UP1 M��ǉ n��\)�Pץ�(��V��l��6xbӠ}�(<YZ�T�o�<uxI���?��5q{��Y���;͕����U�o��6l� 0"&.�;���� t5t�(�9��,�k�8�)�����61�D��-k\�֯�d#���	S'�C��	�R�`�!�w]D?���s��_XCj�^�w�Ⱦ�7����NL' BZ��|.����0�;tz� ��E�E&:@T��K�\����

� L��^�oК�2>[i��>$�>����\��4P��}_sG��}9u�gO�[�	m�>W�Ϸ�C����~(6|=�s��uh���]�.�9��!V�z���t�g�r2V�/'�d�ƶ��RE��H�!�]�^�����������ۢ���HߢZ���c-��wW�޲w�ؚ.�#��K���$��i��x!�^u)�/-]OZ�l�7�����u�`�p�}�>��#��1�U[��vP`����8�3"������j)ތ�d�:j �k{U�R�s��l4:�D���Wh:�wM�~|��*�v�����+
ϗO�w/6n�՗� J�:OYR�2�Z�s�.��V8 ��.�(�Cn%�qio��AZܽ_R���^��hC�P�RN��{S�O!����d��{Y�QO�5g��(̪��w�5e�����f�vl/�Lw���d*U��	`�(R|EX�^�5Bq�f��C� ��1�^�ʾH>��䏹�$�Q��E1��w�Fo��ILD��N�l/Z�����h���\��mOd�^���xV�\Uȟkv[���[1������Ufl��GT�T�y�YƏ= q��)���[:i;�/���뉲�d��Q��l�~�;���Fx�O��j�
S	�3���!�ɳD�<���;w�K�j��z�~L�Tݩ�� =�6�<��!k�J�t{댎�G�X^��������Ͳ1WҮ7>]f�PXƘ��������s1s�A1�=�27�(\�L.�sQ7���L�8_���(��f���z�R��q��7�d� ,��Q6b4FAn��m��D�x�*PD�M�B5�?�[{{��/>�q=Ue?6�'R��p���~�D��ˉ�]��a���6���+�9M2 ��S�p�h����+)Fv�6J�
�z��ױx��󛐨���uyoo�N�V��Y���-F�Yz�ʐ�ah�Q��MV�9N6�py�`GH�~l�{�kf�1���8.��h�Ú�W|t*�#A�W���o�aT�i��\F��O�H��,[F�ׂ
<1����$�h�;m���D��nx�9�bb��}h�,
#]�1�c_t\����.f��_M�0�G%�Y��_��oɓ��tP��6|�}�usx"��4ռ�t�㇖}���{���~�'�Y�$1fVv5F��|� �߭�(Mڪ��L��l^ � Z�'k1�̽��S��r�)=���
Xu�u��^�R��T���ϠP��j��.�1W MCP���\�7�!3'�Y0����˦o�Y0QU���?��蓽�����ɠ��8�F�(Q���)��:��pס؁�:�9����T��v�����O�h�h�����M�����������Gi�����f69jE��ӛ��P��f������7F5͵�7I�\���