XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����b�sPs7['0Z���\M101�U��o`<V07�T]�5�?�26�J�8�g��j|
�ʻ:<wy#=�{UP��מ�<tim��g��ח&�����q��K>S��i��2 �����n��n�����i5����f"��A�8R��c6q�t�;}r�Ԧ��|�S�p��)
�zq�7�~��'���ލ)��@8U��;pRkb�}�B���(�b�6Sm�;{�Һ��mWu�k�6�����v?��H�`M��TE$�L?�,�&AB|Q����Y3�$Ue��4�c�T��NܽW�]��D��Yn�1��[�:ܝ+50z��7��c�~�M�Ans�!*i����^!���@px�4��{w��W��qyG�`�+��X
�דrȦ���@�%f"�F�E��q`"���#�4��w�@��u2pG��#�-w�8�Hdz*�DӹpzE��ϙ1��S�V������y�P÷�V�W��e�:�����V��Tn`m)(�G��0�^��1�rE�G�-[�(5���ȝ~v�j�݂2��!u��s�6vL��H�J�~L:f�Щk�{=�%r�~\�g�T�nJ���x�s�F�E�����n�x$f^��3�}��9�xQ:G�EB����i��.�g��󆆄���L1�ڲ����t�D���<:��\n`�]���^�o;���@IBU/tBsb�D/8�g	�!<��M�����p����gH�I��>�XlxVHYEB     82a     300���n�1����h-��Xa(ڧ���������ȧ��eO�m�b�����:�.}�f�Y�/���Sݙ֖���
�P��"����qt��-��X
4�5`3���y�6�
�0�p��I:[��������MR�����1�P��M5�_W��<$je���I�~E�V*e��.�%$12y�K#93���*yS��g���ZM��_t����;�)&P	�7�n��]t;���sv*؋���W��C���l��\�κ������O0�����x7u�5W\MQ���e�)9�j˞'�G��R7���SG_*�}t���]'�=��v{��H�2����z�3�&�w�V�����č�`}�췥p9����#�>):�G)#J8rB{�M$M���Dxw|"7��Ѩ'}R%V�5QO/�t^�'�S�>r�{��d�6E~� �{� M�#�b;봂����g�]�Hw�<�KM��䤘0/[,��m���QoY�L���;�T���к-�a���@�Ax�cr#�<��Yh�Aʛ"�y��c���HqN,��#���ŉm�Ш~����;f���攜�Z\��1���_�ԶǺ*�E�����V9Zi��^�KVnQ���F8�P%gp_��W�;	މc2V�e�"�ך0j�	*�'?�+&�˪}�����=D���=G���>ּ�r����E���B�C��[�Ecb	O�V�����yd��N�s�����sc#htk�Z�%h��ԃ}����
Ҿը/p1^<