XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Ckxwkv�1��=���Y��G%�������r�3��P֛��k(�ց�r��>!�[2O0R�3��U�w��B���&��D3%ͭ�=�2R�z����Y��5[h�n8�LϩrA$f2�#�m��[����[��#x��Ho��6H���c�������!q�#L������&�f��4z4^:O�{����`�q��7πn%��<��~0�j�q�c�ܯ��<�aG�c1����<� P�-��=���>�.k[���׾hĒFYK�i��z�pU&�fM
�:�&.	��`�BZę/�<�Ʃ]���ʀ�-R��9\��r�_X�o~��+lQ���
����7w��|���yjyAd��$�[�(Щ��;�a�U��� 7��I��-��������lu�����:\G�m9�
깠.�S����>1����S���k
�Cr�+��ʜi��Z��S��̗I��u�9(	5�S���Y�njo@
/u�� �j~F[0h@��HEq9�3"3;Fk?l�X�=�kW1�Ƴ�0�n���n��?���GhB�,;��0=�+�r��
j�Q]pu����}����H��_�0�2�*Ъ��9�ʗ$��Q�Wܩ':��k��^ �J �ɣh�
$��^��Zk9�בu���y��PC 1 RK�J�y�ա�6y#�r\��[��6(;�Š�]�}H�A}��������i�Lѐ7�H5p@2��i��q-m?"D�!�7h!�����XlxVHYEB    6fd8     c30�:ܥaϲy������3�O���3��j�C18�賳�?-Ys��7v;qz��"#�^��i���<|��G���]��7h �ЧC�9?qBb���MP?��=ۓ�.^ 0�or�1��� w#v�8y#>e/�]��- ��]�k ͵��r �hӜ�,&6n�C����:�A,����HQ8
y��?�5ܔ��,5���dTM��s�ƔEI��E�"���E�E�����!>[\a% �Ƭb�F(����mɔ�q�J�:����5�����Ȑe�2B��Ƌ����u�}����:�q�m+����T���&_��j�Wɩq� �9h����#�Ш��,�k:��a�t��o��E��=���jLf�%�:ioo��k��=�/�x���?;�&��&Z]��TO�@�}x	_&k���cT9J�M2�ذ�k�J[,��5��O5�k�H��6����/�[�4i�k�86$38��m�_R6Z1�դ��^�����M#�������
�}}ZϤ��=��Q����>c�KN���tӢ�V�m\)0�<'񑋥 {�H{��7�(�@�ē,�q�o�i�1��1�g��r���$�ٸ��T�%Ϻ>֝ő�R�3�Fw�Wo�x#�_�V��	�>�X�)7`���M�+ ��`�� ��r5��D�@�^Ӊڍۯi)��꽉x�
g5�l�?r��������jH�����E�U�d��q�2}�����,�Rg�)��#y?R����JM�/�`q���P��>�B���ה����N#���]������bUCu�����ZZB��C�Z�������wm8f0��n�\����7=��8��b}ط~�Bser�(��q����y-c@�FG��`�o7�A��J ͓��� ͑g:�=��d9Y[-�J\f?6���6r5�o�TL������a¼c�r��k��6���k��f� I��0d�7�u�ݍ�v�D,�]��(��,Ux����,��\:��.�AޙA�$#s�!�|�C�nͷ;<����eX����lsߵ�gnġa�����V�h��'���IA;9 ��?mF�[���c�b{{�����x�;2������NA��׸ɥ��)I���C�:�������= 
3�;M���B�Se���1�p��8�� q؋�W��~�16��Er�%�����O
�%\%��7���@2�$��F*ѼG*j�!.P�<��>�ƙ���3E�B����'�BQ�o����z��{����Z��T'2Fj��ks�.��C�H���ǆ�頟OܡI�n1��M���t�:�����Ȃ}ל�g�7q�o�n�=D�(`�W
��	 6�k�y ��2�4SV�O�]��Ҭ�#����<"�2��O��Kk�T99�*l×�j#"4V����Bi�	&"�|�k�h����|2�է2Ծ�˾���mv��a��
���R$� XŪ��/�?~մ$�Qc?��>#�r��B�c$J[�&j%C�����*�O��\σW�e³�F?O����®�u��yk	s>�C~у�B�ߕJe�W��`������k�IØ���D-G�P4$��m�>q���#���[���q���-Yb���V7��;�"���;��i��)i�U	L7�Q+����J-��6D�(]܇���D�x��g�%���D��g4����lߙ%n���H:H�c�ߩx�귑-@�TXivun5T�B�l��p�3�e3��)	t̄w����{����ی������:�&ԡK(k�g�$[R`�ծ��Sfv�q#�ǆ��qw~f�':�v�CN^�M�آ[�o��sC+������y�)Q� kSe�(��7p8G�̕�f(磹���o��B�� ��!?&�v��
�^Jk������y��A��������!���e�=ȁ���19ޚ��N����y�l�%�H]K{�i���՘ΰ�κwD�N	�fKĴ�:|a�x�nPL;g�[arP�8*6����p*���g�\���R5fL}�g4.�
�)�tй�C���حZ�&���	�8��q�Dx�]p������F[���=P!��{ĸ81ȅ�EFH:L�cz�#{���ܛ[��އ�C_=ZSIw�A~=UmC/[f����Ƕ4�_�W`4���0��d��2YEs��~���c��f�D�b��+�:�����m�ԩ^/�6F>��$ǫ�߆E@�^y��&������d�7�ɘ�UFX�m4GlSh�+�4B�3�����Bqc ���1���I9�v��r������[�vǀm�"m��$����RVI��Bj?ǩ�؟���.\�$�Q�AW�@��� ���� �m�S����M� ��6Y��f3{W]��uk��=Bf:���-e�R�����^׾������2�)I7`D=�t����&�S���&���$�b�G8��WN�N��Dyuk����&~�=�<|
o��гagA��|�q���'%�or=���w��+t{��j��^�Rn�36�>��<�~n��H�)���١��R	�۟i�k�	d��ZT��j�Șg�3���]�XB�P�Ǽ8�'�Ge2�R�x.p�p�h���.�\��u�Gr��?��:��b`	4FT`����<�>��5T�^�����t��p�ZЁS?oW>f_��^]�FZ�_H�ܦ]�m�Oo��!B��2�׍���|�qے�0ٳ�v]U���, ��7)7���LI[^2��0~�'#�d⢨��������1�J�ր �tf��U�fv����;�ĺ��?2}����3�|LI�+"��Ch���:pl̽)�C�dlgjN�U69m9�O;�0�a�QD�UYN'�ɤ�&��Eɯ^h%�
��3K�;͒}-ѕ�\1�:^�� Ub���~w�>�
��H$�;D���)s��Yw�/��������[���S?�z�����h��Y�% �獮�}0��r e�:��;�s��Z������?76�3�v���{����\�W�v2�X�],-�&|����T��9I����Cec,R(QMKگ�ۃi��}��T_�jJd��".:ڟN<�O�n�