XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����ґ yğK;�e�\%O1%�P���b����4;�#�d��?���GI�D��8��a�5u�o��k�a�dl�),H�=�� �cC�c�Z���$8qo�R��j�È1����J�C�J���=�̳Ѽ����;�|BL��z��x�b��m�R�GRj!S3b�������(�/9 �	kS����f��<���Sx�1��� #|���;�&Tհ`!0�)x���eɹl�״Ŭ�h ��ס��lpw�����r�)x�������>�L�/1�-���g�Z�ã�PI��&�H������q�� �Xk�V_I�J5��'/�N����U�����b���v��J�.<���4��̤�D;s��7��6	���N`�K�K5�������>��5�}��ɍ�'EA�ufF�Z/c^,�"�gv�'��B3y���t��%���t#KaL��ӫ��mT��n��$�Q��]Z'��F���t�r1=L#���G�NT1����fL��V���6I�D7��|<^s8��'g��D��3��3�)���Ʋ8`{׫��q7�\�~��~)�`���9��X��{@�m���Df��~>�)P�A�� ������3&S�,�)�ܐ�Y�����2�s�i�5ќ�����l��c�~��)�9�'r�s��1(A��p���E<�|L5{�LX�Ja�`�+��_k�Q�Z۪=�Ƒ^��&;�[����z�vw^d��Z���<�R~�s�ЈyM�XlxVHYEB    10b5     410x�|V�̶���N��y2>4,.���zR;S��f�6��)��'��q�鱸�܏���l ���_ ���`j�t��l���:(�~�ڀ�*�6�@�TqVB�I>q2G�)L�|)CB����Pt���ɨ��7Y6.���i�$]w�9��%s�+sC�I��0�,�M�!���AD27��R)
���ʆ���)�sh:�E ��5�X��"Qڻ�	w�K9?��|����J;e~�!e�#rp�>��P�/��X�1ݟ�4��0'��	�Av����v+9��x���I\�B BD8~lm���;j���)*5�}0��_�޳MA_0���h�Əg������6>���G��r��)����Ri��>+�t0@���1�t� S��#�a����n�M�䅿P����mBWY�t���}���8���|��@i^��v�ez���Gz[�H__K�[�Q���f�[a%��}��6S�*w[e��.�x�بF��T�Ҙ����R�h�#!�!�#�p�� kPR6����b͇�6��-P0i�Q��Wό.�2[�
��ƃ��(�G�B�f�B#�1�Ɇ�5��:��������bp�J��G�w�1M�6���/�aq��Gw+��,���3_��m��������c?j���8�����N�pޮ����a�a}��?ZBxW0FC���PA��JK~�1V֜׌4�[a�C@�Eʠ��[��=���*m�,f^���Pf�p��Ds��p��wt�hw�zpi{����*$��G"{�����G�8�Enēd���+y:׿y�P$&�ٰإ�W�(S�Ð.q����r�.�5�IԵ�h�"n���>UZ[�a�.�Lrpb<-��20~��������x)!�km�˩�i&gި��O��ԍR��|�y��5�3e<���NM�?�g��o�r��[�U�ڼĥɷ�^7^w�lJ���k�F��A΍�ŀ��,	4!�Vi��"8�w\z�A�GI��D�Eϵ"I���qP�4Ɵ����!�`K