XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��8]�Je��K�7Z�)�׮U0��]���+�:�=F^X���k�ө�.y�p�<1�Nɕ}���Y	�M
����p��~�������Yf0��X7*�[�U���/9f���ĘĻ�|fÛ�'w��k��Y��kY����7����#4(9a]z^�} �y���v���zW�L���ا�ʓ�q����|����\��ov|c]��v0ǜ��̠~�/�mJ%7���&x�~��{+:��;�u��p4T�)�e�'���wW;��S�<��h�=���IY^�t�zB�t���
ʛ��*���F䗈˗���w�C��o���KBE�)I�EӍY�_��v�k3�2��E��fm�w�p�.E�B����N���н�6"����-p��>|X����`���#T��@f�W�j�t�{������ �xm2M��XS�Fɧ��J��Y@��,��?tS3��P5Q"��k�h�m��:�Fd��#ƭ=U��B�_hg=́D��d�

9h��C�A�e�־�W���ۏ���pw3��6"8�_�>Tc$�X��0�.~f{\Z��Oʯg���Q���tn����v�E��އ�������&��u%�<�U^�c��	���G;+`�$3$�bR�2�tZz�	x�����_���
-�+���p���R"ɢtI�)��}~b�4q��VBm�����ڧ� +��8ssjsOű��iʦ��g����|�z
bǤ(���J�;|.6� ��XlxVHYEB    1cf5     790�un�f<�@Xl�����	sj	�U�sG�S�x�̍n��kh�X�\}z˸&���T^t�8���'��h�!�μ�{�{��4���K����R(
m&Aóe_;�$tPL
���@�| Prx�3�֚ͦ�S�)43�!�ۧ\�`�����Q����Q���P�i=!7c}�p]�����_�J�.d����+�1jF��{���`	`����W�91)k�~����c��B�D�C<xa�j[�,�7��ML'M11C���o���2Ұ�o���J���@��>��O*�m�x��d�=��Ջ��~"��{�7D� ֟9�� ��V�tD��&���q)�����C� ���ow�T �E�FT𻱔��_p�l��PӃr�"�h����1ʤ^�E�oLG�	O"�Φ��,���iF�C�盌%�k�\Q�m�je�w⪵FQ�yP���x|���qNb��d� W�������@��\(֡e���9��2\j���ykn�E�և>�؀�o�P��|�0j��?�΄�j�F}Zk�:�]��c:��5C,�#��C��(pH��:�;�+6i�( ���N�U����	_�?�P/�f��, l�$IcLF��:b�вX9�|P߹��.w����W9$X�����l��d����տ�7 I�c�����f�HF�Ą#����vz���8����W(Z4�-2�1Y/��7��Y	�pN��^��:kdl
�
���s�/k����H��ѻ�t�5�CĊ��6��|k�9�Y6%߅K�IX��}e�i_�M�C6�ڻ��F4�������1�di���ANCک�j�Bx*+��25<~���E�p��|��}�^}����!���{�=/~���8��ǽ4tZ�����y�M^�h�9�$Wbǡ�õ��$@v���*��4����M,\W��b����]�S�+�D�S��/���gV�f-�x��D�*-~U�9�,��@��`���WQ�^E����GU�����w�{��т�sۘ�Ă�d?]����2�R-��)�c�i�!�a���90�&�)�o�b�b�%j� ���?�݉l��D�<]���u�l�n�8���M�@Hk/�(i;8�nV~�
����F�2f���f�!O�sP��=2BszӅf��a�����hx�G��ә���x��K������M\�����J�1���3���
�N���^Q�|v���.���:^=�}XO�� A'?H��`o$�S������8����_�,y,0D��)m��&��L���b8(pIJ��� _�)��
E���`�X@@���b ���R8��FY�P.Sh�
��o�{3�����}�! ��f�(,D�<��`7���n2�'3R6\��|<�r����,�$$ۛ����A}�We����OuVZdʏʨ����|�FJ��	�
��w�n_9a��j�����pK/gr�S��[����\���ũpC2�=�|
p�9��o�&�����\�^D�t_VyS�9M�>��� ��T�=z5	����nN+�$bc����{�5�?��A�F�ĜM�5Ux�FhN�V]�z�����Z���XF�=�{�]�Oq� ���o�%�q?�t�^_�:��C��eЁb<�b��Ӯ��)G2Y��.i`7A뉝�p��Q�l4���Y6;�Q�JY��ֱ3�j���0�-r�N���?�oJ2c�����-]]�����p��;�+�1��k�*���÷h����:y��m9
#���C���1$d���ツ`j�:3�����3�ݴ�J<��6)G�և���d"�D�3@���>�� ��c�Ţ����?伻(��~��eĤE���S�w~�/�o��N�c�?��Ne6<���F�Q��+�!��.��DY_4Ɩ�M