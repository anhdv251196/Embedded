XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��9�o��v�6����ᗙ�EC�l�����q��<4$Lp���6n��������of�v����˧J�/m�N:]IcU�6M9���M��YV���b�>����?�J�)��sV|�<�T��Щ< ���`d��hz{(�K��׍��W���Ŀ���V����T�<?��݁;]�F�#'�9Yj nTC�q�1K�@;kH�������Z�N��or�o�;�Yi�����>���DkuI�?#��b��ޤe2M<�l@�KI�XxTS���-�޹��Q,��j��K���M �����p/L�Zk�sb�h7ڱʊ�v)��7� QS` �1��ƶ79GW�B����1/N�g���%Șϒ�܀1���Fj;u��5SX3(_	���SWη�
��)!�&����fHO�Zi�( -i�kL\�(�Y�h�����%!ř�d��_>�o�{��jZ�jpK(�7��#��
3ǥ-_FA����l�g`H%xu��ت�*+i7e<9]9��yU5��e��2�JlON�l���$��$"B	��VΦ��mD.��~7�蛍�C
�[a����A���14�����0jY�͈V�F���jؠ����!��gL�ȭ2ድa-;��(�J͸H�K=�mP-����u����گ�7��}r��%P�����j��	pq~<)(�\O��X��MfhG i�W39`�d�P1��M�]`��o�b����i�V��6.�ˉ�pQ��&�f/XlxVHYEB     6c5     300�d)�a���t[)u���ۊ�=�܆!:�Q�ĩo?Y,�|2�o%|��RJzK8�o�Ε���F�JӦ��>gg�'\,i�Gs��;=�j�����y4��8�s�Un����I�J{1:O�.>w�BkP��f.F�S�=��4*�� ���E3[v�M?�6vNvcN�3�.b:wK#��SF�����o:/�J��7}^��-�u�P���]j*[wֺ��Q�V��o�ŹQo���Q�Z^�d�3zV���2��3�j=I�IM�m����H��۟�o�T$]�!T�l)w[�rҲܠ�d�RT2�4�P+3�j�3U^�������x���R�=f �*���q�Ϲ�I���֠,���Uj���*���N����iB���m3��q#��Ј�(��i��J�d�pNm}�v��V�]��K6�U��l[��bkh�9�Y.H:N�lZLR=#3_�,�.Y"�KU=#Bf��\���J�7��r����rP� 5��wȜ�0�'g5��YT�G�4pM��q @��Ȝ���#�͘�O��wȫ��+=�3e������B�?�������\jy}wR��9�+���&����Ds�|��e�v�zsm��]SRޡ�leEp/���o�i{��	1�Hc�44�+��o�Պ�J�����qSe��9܋�e���(U3Ϣ{Ef�:�Q��~]��g��<��s�X�'O!���X!�q!+�aNT���y/x�|
