XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���A�x�Ӥ�ĺd����=�����ș���f��K��ʥ�K��Uu|���G�܇M���i!�G�(�J�@\���pCZ��6?%��5e`a�=r;|�'��L݆֙�5>b��^(��ߏ�!=w$dN����	g��N~r���2:�0�4�f!)�X�=;it���`�=Pa�M�Ⱥ�O�Iu�gپ�C��72N�Q!�fS��xFl��d�,t<�|�~usH�h{~6`6��ޮ�,��z�[ʆ�.Bog���c���f���̸!S0�(t�A�K3�[��a$Y�6ܙ:]���}�["=pr	>,�UdI_��(�d�"��p�j��<�s�ڿ(+;���/��nͳ�zkI_�烟���������E简\r���q˽�jX>h��\K�Ǩ+O��_0�)����"�͂���<X�,?5�D��C�K�
m�!��ѕh�(bBW��=��J��W<�8���x�"���)�(L����^(�lP��R!�B�$ [^��޶��Au�c��˭~Ҙ�.X��ꚽq"r�*��5y�"jnYyV��^/�&�܌*	�Kl:s�b�5v��R6�.z!��ih߶�A�T:����1��YF�������`���:�`+\c���Bv�J�#u2�%��[�+,vUڈc��~O�:;f���5�{�B�5(�e�p��ii�η3�TU-T�CB-�^Bu�/*��6=�k�F")r-l���M%L�sC�a��bn�E���`%�C5����RXlxVHYEB    1cf6     790����$����q�׮�p��؞T�OfM��p�_�8��z�}}~̀�O�0W�_���N�|�Ӽ���a<��E
l�J�i�C/�'x�:��XBK��w�΍L�WOp)R�Q�a��۴үU�����\�Rg�֟��d�#S臔���'2[�h��7��^6�,$0A����rY�OJFl�Ψ�^;�����"��Z��l-`W<ވ�����]Y�������0p�C"��O/��A;D���A� 5�4�yh�]VDJ����}Q�7��%u]��M�k��Q���<�ex�pA����X���W����wW�����LtƇ4Bm�����]Gģh����!� 9������1�ҧF�-�y�0|�-Wȱ�3�yL|Ǭ𦖶�JJ��K_��k/EƙV<qfE�1魐��{�Q�5���Np�6W��X�364�G�<�`�������G{��+�P�i���B�CZ�$�����ܼ�ȨS�l��V��/bq��bWϼ�#���F���e�X^���_'o.hi�$�8 W��.��Wr�q�yT{e�������W�niI��9 ��VWO�gI;	-8M�1���:��U�*���'�B7׉%2Έ�L�zN�^�鮰{���`% ���"�kǃm.��"q�\��&��2�'لn���5=`uf���G�{�q`i~�ѡ�)�g3�0�K��@E® t�A����	�Oloɒ���6�sʫy�Y6��+�0�OH9��O1St��v�P5�����ao?�S����5y5~���L�vX�����J�?��X��������ɐr�Z�i���/�M�if!����
�Y��G����T9�>�] ��$��
*�Ѕ�E�e�-*uˠr�	��NG�9�u�H��Jo+�_t���fK����E��:��lo^d��R���4���6P�|W���C���Q���V���s�t�:a��_GvP��^(����r�M(L�m��=�[�$1ĕxQC�zFrb�N���1n5{�ҲjN���]nf��QÕ��k��,sA����.��dݟ�c�>����?�ξ@�~c�5p��[$8v�
!���0��{�2��_����{�Ȩq����P��鉡����9<�G&�{���Cl>n�T�%=(�+��\j���ǨM�.W9'�'�f*ȯ�Oz/՚��1C4j4�̑�/�~嚌C�4F�"K�;/����y�|\{��6�L���:�-�z��M���K��u�Hx�tI������;���g9�!�w4�;9iv-y���1S�7Ga�� :ʨ8�9�L���|��>{d��p\$�B�ѮB۟�KM#[�8�`J�^�b);�"�����5s�z��cx�tDE���QT\̀i&um��D�e�������_�����d@��f���j�b+hs�����0�(Êȇ!�������V�#f6�<��2�q��N�����pŧ��Τӱ�t��1�k��%=��I]_��<6��b��A��1�R-�Ba��6�b�s���^�EtsW)2[�r5�|��[Ձ��Zt��3�O���;�h�B����K�h���t�1:�u�ޙ�z�#�f�K'�k@�%���2�b�@�#�o�[xP��3>�-V}���0���P��8��EW�~�b�����.,����m�R�S�?"�Gݵ�K��>rr�j��k�jo'M�4�3
]��u1�}z*���r�4&�?�&����k�G!GcOGNށ����S<f!!�i��< �{ʴj�	}�D�n!9����8�/w<��
.7�������T,c\3�-����[ ��*� T��繁��N�1ۇ�TY�gx$v�D�
�eH s�O�dU�,��M</ai!�H���j�w���)��Zx