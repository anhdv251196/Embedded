XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��P�2<�,rgW�w�^�T۩x��7b� (f�oyL�)F7� :J|���\�}���H�c�WOA�J���>�� �p,�2��������&$ާؕ���a�j�����b���D�����Nˮ��т<�	e��S�.���b^�)V�����T�G��E�Dt������9�&�젟o��E���ן���<j[�0��UY=�'oc��h#�8�.��1��_mA�5?�Q�+��4��l�d�GL����Y ��Z�a�pI�W�aSg��=���x�H# �ӿ6B��M�6I��b&6\}NK��Z#��&��b�Ӻ5��V�X]��yZ�fE��:������z��K��SЁ�Ev��
��k���i��Q0X��=��D��K%�BI�b�V�6R1L/èp��K/�!F��-,����L���a�g��!�jQ�N~��o�1�g��iP2cF���7��w��UAW�Wa}�D־Jt{�1�j���[��C�	�����S�$	�Hx�E�I*�k*{|~��`\���L�>��&�˾?R\��+@�ib�U�W�Q~*s���G�滤l M#�zHʔ�	ax��-$��)d���s�C��r2$_��g\���u֨JH��A���a�Y�*ɋ̵p�|�Kp��Y	�΅'I��,�����H��6,�P!�ia������I��nO߸q�����L5}z��C�0�*fj�:�˱l�J���URQ�N��u��[re�x{��('�͍y��XlxVHYEB     a3a     370�R��<�p�=�
h^���Р��+�#&�8"7Ftu�a�$�_�gXR�
�Q�I����|��0�2���důZ���;o9��ߍ��C%��yz�'FF�&E6���j�d*�9�7p����k�E�*s ԰���T���H����{
��3$?^�vUX�s6Ä�"
����v$O!=B/y$'+�hr��,�K&7�{l3+
��O�x����l���>��gO?#�_���y�t��^�y�$��9R�u�P�T���.�HP�`-���#�ڕB�� _C�P<8��QI1b�h_�:%�D�.8xtRyd�G4��xk0�K��-]�N�	v.�U����M��a)�軀��ٽ�%�/;����D�}��Ѭ�0�\�7.]dR�m�Ur�v=鄕��Jc����,W)� ���r7ނ^X��<���)�ʠ�}l�i��Pz�I��Ԩ��Lc"M�v��"�)!Uq}�ӊ���8x������~9-]���H�!s=$�ʑ| ��R����`��Ekj
�ēb�f��Tw���rb�g��i|����̃�W��On5α:}i��$����UUO��+W�Hix�%0	�#�>	�Q�
掫edTL��z�GI1fC�]����fdr�4Rw]��n?�@Ǿ�VWZ��RZ,
�b���W����."t�h#\6�UET�'�Zv����s��j�����Yܵ������[����U^��+����ò�Cχ��t' ɺ�A��/�2�O��o!!:��ȭ��H���te�6�
$��9�VP�\���u�E� ᣐS���d]c
nR���5��T���R���@:ip'� �fF�v�w�R���V��R����ǝ��