XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��'�SJ3�����S\���_̱��3MJa��96F�w���a{&8�`7�c��9���)(��^sp=�g���1��s�Xf����?<o�� ����D�!Fs����S���/t��W]���;�Pm�y�o�4g��{Q0������8Ո�z��ANºʶw�L̐ս�jX������3:q�­>p����~��pG(v�X͊V���[��Y���o{S������)m��l�U�e>�C6R:��t��h����m*�<���Ef ���^�ܴ�i�Xo�	Ix�lS����u��9(~Q�ڡ���I_���Т��o�)�U�!��� 9TC^�]�ƞRxn � "�8j�=�Nab�����F.+IDz��b��.�̀9��W���-�nŔ3�8���X���z��eIJбoy����Ǐ��v�'���!���bWi��?���������2��Ӫ��'�*-����7@o���/Cm�!�xW��$�� z�:�.ϟ�)�b3�ȩ/��?�˵���~�#�oc��hB#:�Gx��kЏ��r��E�t֗!�%�  �k��9U<2���򯉻��´�otC�7�:}��
l�C$�*{��:�9��n?l;���B�G^+N	\��z�n��E�#Р)+v��n�]��2�Ė��$���a��C��P	XY��)��B�}����W�'0�S55�����h֍��E�Z�he>ce$���U/pm,�$ü��(�;��XlxVHYEB    3248     930确FrG�@쨬$ ��������e8���HUHP�.ս��/�8�=
l������5�F��G|<�_F��:��{�v)Ls��~�8ao��7�,j��C0�5�	U�e0%�4�De�\�g�"��\�A�aG�h�cz�Q�sU����+�v ���QSE�����zB�a�i��ZY#ԁ}ߩiK�9����ه]�2+�*x�W
�iȹ���=_M�E�����Js�o�E�:�:�<ʛO����a�Yh�9XS{�ovyj��iΊ{�!�?J�/�� p�U�m�w�f)��G��:x)���5}|r��rjR �X$b<���F��j�Vp0zF�+!���e�|d��'P׿-k���I�3�X	�!�]g��
L{;l�4Ĺ�%�jI���6�[��F��W:��u�k7�K?�EFC�R��&d�`�Q��}Pb��ζb�(�~[�l��:&j�G%�@B��b`��~�#��?	ő7����x�gM�R���7N��)�ǟ�sS��a�2���[x����7�@���87SPBxܗD+F�Ve'saT}`ߗ�˜V��Y��C󷁑 j��A�Ԛ}���⌊�7{����&6T����`'a ��$n�栈�]��v�3�w-��L�+�LDKS�Y��
�<eky�23���X�姽T��4j~��n1�g��U�!C��կ@u��ȓd/L��Z�{��9�Œ�^1$���N�im��]LO�U[�D)P��Lb4�@}����z̩ǍV�[�x��g`rY� >���t
��#�D����A�	1�>�3!'p~s<�p�Gt�/ox1��@)��ߊ����)���!&�c:��I����j��GW$D�#iP���-�R%6� uM�<;�&�|0�B���i��x�6G��a�t��ʂ8h�y����L���	��[M�r�o�
�����
��QI�$�D�y6-��(z���X)�R��J���sh���6�T��}kޘ� ΅l�j,�%���A%�|�S,�02�`r���R;us���L�oQ_���rpC���;��'n��VqW�����l8��E�$�6f�T-ߓ�}��T�"��E��"�K"S�Z�w��|i����.>�a{�?f��5c����"�`4����f�܄H��g�MXq��������ۀء�0
ļ�Cdb `�Ɏ�2�1�{C�s=]*�g�+ݖ��Ӌ ���oۙo.�-f����y�G�ųNp�C�gh��0nLs�t;��fϡr�˜0��qg�~��bk�iW���Ӑqb�	�qNIǿ������)ͬ���Rmn�����|��u�ǎV����o*`�I������2В�.���g�?�S����<H��U�j��}Q ������}N�̨7a�~��"]!/�p����g+��/�D�ֆs��0�F�E����h�x��x�j�PV��է�GP��HҠ�.^�;�5��F�\5�`V؟��K'uBs[��Ҁ`� ������2�F]�W�3Hϸ�1��ݴ���h��u�7����Ob�k�N��qP0����P$�#��y���\IP��
�}�O�@;��#��a���$�.�KE���>���	m�?h3p%�.�q�vB���uI���|�����$��(_;�3M�T�����1�`p���r��}�J'����(�i
Vc|,=��.�K��(�f��IU蛝{r�ToòO����'�O���Ꮣ�+ʂի7N_<fz��gw����(�9j<"�I�V���6��6֌4Fz�?�^v�z�b_�C��x����Q���덑��w5��`��
 sB��~b����-��|.�5m[}�ģ�Sɪ5j�=/v� �)�u�����J�N_��|�ϓ#����55��
��Fw�ɹ�=O�lD���{d7�>8�(�����U �r|U<f�Ut:��u͆a�)rɡm!��}��(��0*�khI����B��*X�]�c�����b����ze���=���̿��:88�?��
nO����*Ӻ���V�����⣉CVP9�-T[���U�P4�j�K�ɐ�l�wuq�U���n�4���;)?X����ʂD���mV��� ��������T6?��Q�����z����z1	襈t��Q�\7\�N��,D7�mC�`!S� ��Z�Tu�E��?{�R�&б��Z��m�3����Zx�����d��E�P.h~�� s<l��M^��o&���Yض���\(�����O�DI]�DI��h��}��`��M5-��`��gV�����G�|�Ń��
˦��B���