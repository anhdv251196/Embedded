XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��T�"i�s�=Ǵ@g��6��z��YJ�q9�n�qh7� kj¼W���8^3��l�b��g�oo�4�S� )��U��j��<�w�����׎eז,�����W�~qβg��~���|�]�%S0��X�-_��a7�JN��3�1$�9%���'hc����=VU J�=7P�_��PvO��7�*���8�#S�I��|�����?������줶V�N��|�DB义�՘�Q��&����@�pi�����[I�=��U(:�+Ϙ��VP�̴��p��ҋGp	���ـ�J�Z���[=�V�<zS��`�T�+��=�w��_]M��7P��Ѩ��h_�a�x^�_$f�+��5B#ۤ�VL~�t���UNDe�����4���p
͡�*-=<���i���U~=G������+M�3��J��@_�i?�v&����ܖ4Y ��7{~��[A���(��T�ޙ��?�M@�'���Ƶ�*��!9��/�X�\mt[��[0����ZL:[�e̲ˆ��\4�=S��*���'YrE/�o��כ>�Ȕ|��R�:<��[��}yי�#���� T>��JsY:�}>�4L(�3q7i�	�~
�Ʒ4�o��9�(fm����yp#�棟5!uy�M��W��N���aG���?4��̬^�p.KBm�g��6D9:��yv��ڟ~
��xҔ:���s���T�R�*���i�m�X@L��:]H^9�x�BB�sOG�,�ĳ$����
8�XlxVHYEB    11e4     520�b�x�N��)�l�x���2y�T�,� L^��Ѳ@������ִ������H�tҶrF�����E�C�e��jYJ��>L�߯�q���Zf;�1�D*�� �ӀUg�ؘd�,)+/ƭG�����r���WǬy�zc�Px��	(%>p�6�o^����/
ޱf�ܷ!�sV� �=/��zFg�R�|��dD0,)��7ױ@��ɥ�WK3�EϜ��h��?�E�� �pE�bv"�g�H��}�GC��%s������nK��F�S�t���-�k�`�qom.�\�Ӳ�Y�#!n�	Ԩ�@a�..�5��;ay$��x=Zy{��ǱhBR���o��H�Ԫ41k2���r�ģ� �8ў��i��%� gM4 �c�������z���<��r�`��7}�~��*�F]V�`UT�Sgb�D���_$w��!�MXC����A&:��*�r]#v��e�iMJe�f��l�0d{�Ք"���Z�˃gߣT�Q�Z���N��1���ؐoI�Ʊ�Kv�������Y�&�Βqaݕ���6��m@!�u�|?wU�6X�O� @Q��H}�VA��c �<kP?h}Up��Ĕ�n�d��YmHQs�7�~�Q�0è�@1���s�z�r��v-�V�S߂t_�t�l�����|���
���@��sC�֚4Wlz��"u��Z�c:��#y��K��>��sZK��j��.�V Y[9�2��ʍC��D��!}沈$�y�l���l�D�zEC+���v}@��F�&��2���3�
ބ9�Пo]Հ��3� q���2ч�wC�XO�U��p��A�
g+˝���ށ��&����	ʹ��5J[b�O�n+��Rx	����[`j|��X�G���k ��,�d"�NO��dWC�5d�2����T���d$�9�N��6u�O��xc�8
rC]��v��*\h|�����.����L�o��\�V�	������'\6&R��|��l����O#o�g �W�6��}N�اx�	�-[�Rw1�
�ģS�(F+���������EA�#�>��
f��rTèl()��
�y#zg槒�hе=?�qv+��LX�ga<8��.�UY�� ���ꚷ�P�GFҫ6��!=k�#ى�}{q-wk�:���E�.�܂N��Pݢ�9ڧz'�	H�_%��g�A���ݙP
��3�Z�l�.4���Jƍ���ϤOh��Y-Kk͞+�^a��A�Ԕ<�2���[x�P:���?��#�k�#|�t��,�I�17�