XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���\8����]��B�G��1MU9���U�{�#B�Q����I.�<y%Dwt��v;`�x�������HD�Z��o��O���T�驪P��ڻґ�E@d 9BF��{��eP��^p�B�aЫ��_��t�����rX��/E� �(���(���ƁBv�U�5^(p*�Eq	3�U� ���)A����a�Q��`t@+d��� 4�	���]M��欖_�s�fP�����\��e�:~�>�� ՚m�9'ٗ�}��A��9���yC��=X��'c�+�.1�nC��?j���m~��.Bcb���S(�b1���W����T	0P��������k�DVʓ���$	�n.X]��<ZC.�R�q�ɭe�y�S�*jRf����;g�
3a����p��y�А������oU��h���5x��6@V�d�����9p|onQA���de��=�@���ϱ��WZkj3&�n�WO�25R�+�3������Dq�3�`�Vn�e�7��2G���Jmn�D{oNyT=h�'d=h�M�L4E�ߘ9^�}Te�;В�Pد���L�x�����΄a��3�HMC��K�bC}�[]��a���z�.��ȹP<6��=��:/�� �y���2�e��k�:�k_��	�)��e:��k&�Z�d����#��?���o��ldkcW�i&������F�+^Zns�-�hؖ_�[���qY�����MR8l�3�uae]9��q�#4XlxVHYEB     7d5     300�;��U�d�>�f\Yq	����o����k���m����ɳ���w�V��0��Lˍ�yϜ��<�{4��w�s5�\���"�b�xߪ��E��WA�tf�4��2��<�fCt7^����i��y�n#��T�K��o���i��D��f�ZPiB���=��tZ��Y)e:���`�l�8aŗ��?�0��x�@�Etp�cS�������4��.��6+WL�n�:�#�@���i{NtLH�;��h�]��}��|��̉M�B'���;�D\������^���6� Qĭ4R>������Y���讏m�7��^`u~��B��:�����56��*��+ۚG]47z�a_�WBo=u�]��3r2��z`q����a��bE\,�d0I�&͡�aU�]�����'�����+�8�#�Bd�tQ�Wu�\c�^*4�/D��y동UE+V�7�E��玝��b~�q�`�P!(Z���a��3�\MN#~ŋb��`�<�X`���3���UYGC}��#HL�[�N�VU���-L·�&x��a�^�9̞S����\��N����~
��_�Eו�?Tr}�d�&�uϕ)l�m�W��$�"!R��rrj��Ҏ�D}�A�E�.'5�lW4#�.6�El�zn�R�og�]��$��}�&l�@���J$��N	�ܔ��B�c��l�zX�ʾ�£S'���C������f�F��/�t42RT��V������ �of��cjN��v�)�)