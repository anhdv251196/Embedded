XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���ci���ܿ%f���aI�9" ��ݎ}>QEvM@dk���B!�w"���/��1Z���bt�v!�U��Np���Me�{0�`��L�%�#�,;��،��p@��+2��ŭ�>Q�IK��Y���XN�������o���	^I��r�ǽKė���������bIw�C���	�Z9�?�ջ(أ_��/�&AW�<q�n�#(�<��D�S[��DG���eϘ����[iL5/�py�����
�ց��.Q	�"��%���#�'G$H�3���������Ft���Z�0��L3/��
�|C �^���+=C�p�P��1׋�-��]�a�ou��/�y���CZ[$��$�W�V#3�t��� J���~V��nHDb��Z�#�Y�<4��[E T�k�f��xeZ�*d��)u�'i�N�>�J�����v}��#�i��e@��=L�q�0�q7��������`WG�3�i�
�ϔ�2Y�Zq���ˎz��
Ԛi�Xc���M���uY�<�ĺ��Բ����N$BV�=@��a�l�U�t1�
&��Òh,���'^��4�zjhg�`���ja�璪B�����<契]"o}�x��"ٖL;r1j��=��*�k���ʂ�L�߿����k2�v	��H�X��}?�-Y����n#�uZ^�Q<@oe�mꄭ/��2upY��\�l�?��N�і�����vP��!-oT��8�×uN��dNs�pc�ƹ�|�MgZK	m�D�XlxVHYEB    152e     580����$��Y�Z22Z^���:���[v�m8>+A������.d�S���������U��3�c_94��^S4�)��M�Ywz���1�ǉ�0���׺�7��@vM�`���y�rИ1��g�w��론��&%������NA��0ʜ���},� ��Fx�UNn˂���ƀ���J��EH�I�$�o%樧|���^p��
���ɋ���p��x��v�av�T���l�b(ĝؑc/f�Â�j�_�Q_!N�l��r��b����"���u_�9�0trX����"�>i[�e�Tt�ǆ ������!{��u{CM���cp��U5�c�=$�"�Xx�+��X-xf�)����]�6�)�!��y̯�C���+!/��{"w�G��Ցzo~'��g|7�*��C�Tq��R�hS�KFv���T�B��̼����w���봒�'N��-�hH�fJ��\�zO`t��0S��˜h)T��%V�	?�l��wԽ�����x3d�����o�$�&~|�Ĥ�V�&n'ԯ���yB��2S�J6�(<e�A�Cի�a�EN1|�L��wG�o	�8D�τ͒�5��m�,���PV��L�Ⅿ���Y�i��z�"�ؖ<?�~{!��k�QQdT@ƥ\���'��C�� t�[P��I�H���Ãgc����[���w�̃N�-I�=ki��M �L�`�&J�΃�S�.���LH�B)-#ӗ�ss����5�QM6$���d��6`	J�1Є��mGX�+/���G!�O$׈7}�K8uF�g�-x��/~���֗B�*v�1�0va�]@�yw��� �A�?p;0�Px;��S·1%���I�M�$�?5�}͐�ى�{�8�#N�5�l%$�	�U�U}�|��;�����j&Ca�}Se'Ej��n�f7��t;�R3��`K8�4�J'��펩�&A�pZG��0�B�,M�|р��1H��~�q�2��Л����u���n�i!�\I�/w�`� �dL�á�����4��O��ț.bs&����c���f�����t_Q,g���,��Y�P����b&��P"�����zn!�4
�U�U����J��'�)MϘ�]Ӟ=����U�:@�3�M�� ��6]�$4�	�U��KŬ�X�B'u�'l�.���۱��s�'�M4I��kUX��_�jM���'x�yJŉ3���
ЙzSkT�&������)����,��V��ϕg��g(~�?+R�,��,�ӝ"ZP�i�X�U�4sH�M�p3����l���f��f����ˮnEWn�z�+ TҢ���Q@�Vլ����zT��h
A�|��@2G^}�j"�%�`�{'��A��B|�?p�ܦ���u֋��h��&