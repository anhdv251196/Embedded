XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��9m������!n̕���s�p�.��֜�/�����RTKh����S��o��:N�IVRIG�8?I�|9b6���l/ӝ�U�p���͟�ͣ�&CC�ݧ�%,��o���x�_��!=D�� f����ѐ���	0�*��$T��@��_P�ب"�yĸ@.q
_����2��L#�sc���u����Z��ަի�V{�Ue�vx���K��yc�j~Ԕ����F���P���3��7��06���Hn���AÂ��S)������*����zI1�$BQE<�ޓ��'��)�4r���X�_����;Fv3RB�]h�|o.�]�d)�ﵻ��}���'2��Ȁ����䝢x%�niE�`6G��:M'b�<�4%�����\x/W5��P�����_04�ix:D��caSC��%K}��(>�޾睱07��e4�4�׼:ꤍ���.������[ԘB;��u!��=(5���j��sg���&#�%@g����R<��vv�#�Z��R�O
0F"��K`��Ȕh��7b�������F�%BDݨ�ʈ�i������l�(I@<d�6��3�!@0	9q�<� ����!{T)��>K9�1K�c�D�X8��1�Զ`��_j`��I����J�}��A�Գ2�\I~�X��؞� B��v�`�4n]���3���&y,���|��cT�	�.B���Q42/<�V�e�}뀓���%�w|l�a�^D�E�"�m٧�����`3���q�V���X�XlxVHYEB     ab5     420<�R[��8�M{3�QS��M���ZC/��+��C���U�(SV�.��r�OщZ\��:FU�2��Au!(�!e﩯z�J�D������D�Kv����2U�����%��Z�9	=� �%��tȱO��7{�0i0�]7x�/mu	��k�c"o�tZQy䆷��\S�7���&��# ��&N�LN^��4������X!w�a�iC�{L�����'m�Fr,g�5�o�uV\���yA:xp��=}e8Sd��{��W�W��bN�V)�˷��^��$}�����fH]��
�+��}�8����ܵw\�Y��<�:�><��T�.���/�����O�N���*�AM_��
nP:��|�W H�����a�x2���}~Y�fy��ǦK��Զs��}9q@G{�r;[J��c�j�r:��$��+�B6�Tz���H�����2l���S(���:�w���՞�J�$Ѹ���y&�.�����=�A�yK���<�<��U`�^A����<�l���T�p>h1��"�>}R�T�_eBj���2,j���T�7C�Cd��'q�'��,�u��GL�o�	ϔ1f��µԵl���I��R��c��ƻQ�K��p���(�9u��N��T|ڼJ� C$) QPcԇdfOQ�L�&:�g3n�Oݠ����B��+�HC����y�a���J�����o�W�����!Ol�"C�,��(ZH���8ܯ��L�)p^P��K���shg����K0cU8_��(��`�����?�;�{(�z��s������q�6ޔX�5D�9|7�F��\u��^�b�Bd�kK�'F��c�~X��h�d/�a����s�5x�*��I/�k}N��[MUfJo�0��D�j�?�}�T�jj���|�h%��󉮅V��ULΒ�r8M �d}�%��l�s�
��r�G[a��Tӽ�ńu�vhIu�ȿ��vab{����� ��L�:��h�nb�&����${a��`����~��/��f�v<d0�A