XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������1*������eg�5���V*U/��u��@s Kܙ~��ڳ�&�S|� PǨtZ,V�s= :�rYF\s��ō#gR��O*u�����6�Y��{���r�Q&�3Sk���S��s?�:Fo���u]���2�o�}��e��R�6��F����&d�Ug���f_�陳��2�uka�,����K�a��5�S��YM���u�.E(�O�I�0
�&��f��~�=N���R��ֳ���tL�Q���^�1��n�K*��X����0+�bܡ��0�^^�6ns#���צ$����v�Q��]��3���ׅ��7�Ҭ&��7��A������b1C����z���G��I�}Y���g�.��"M�C�ʹ4̶<�U���{u�%���!�VpA:�I����+.��˖���/@{�_�G�Y�]����;�Q�WT,��Z3��L���8�EҞ<���ǂ�݀%�i&T�Y�S�B�]�mA:ǌ
1K���}�΃?��^�&���U�oW�{�������x�\�Ȍ~���I?�ӆ�R��c3$]n���ۖ��Yiϓ���S�?oe:��wi+�}�����{�	� :�п7��<^L�6 X������?'����u��Y�y�51��Dܰ�.3'�{��*��G�$��:`���bd92��Z���F� 	��.�w��_����QZhM��`���
�����#�{�mq@���@�s�����Q�"���FW=%2
�oW�H�4�m�dS��uXlxVHYEB    1c48     560�zh!���9eD�u</
�́�~�0N*]�5�쫌�B�'�-R�sX�>!iz�w0 ��[�f%�t%�[�M˩@!�d+�ST>Q�Sd�r����	��̰T��ʘ��t����R򍥗�B��2��ތ|�$���H��f zh\BBz��F@�!���<�H�ﺹ���M��<�v� r8��Y�����K��p>Cb �	श&�}�nY��FX_?��h�uoK�2��T��>;��c�vD�D��%+����׷���V%FH	�8�`�c�̷��g&S�����p����wwk@���}���K�ղ��9f\?�6�Z�+`���.�Ρ��ߍ�HHn�����Y;�`_�Yj����i"�t�lm���W�:@N�ߐ���Y�A����	��3�e�D�Uǭͽ~�a�G�4
��mT�`�P��[
�H81�����oi~�w�0a��X!~��N-r�Fr�nk���DA��'���/��~֊@�(��]���t��W�<��։y�-NT�!ww�蹦���L����;�̍%�W,��1߰��3�k�����M�9iF�q��i>楧XUe�9���^r��a� ��e�b=�
u����;i}*�u�
�׊������e�p�W� �Y����4��O�\�,�{ytIL
����$	$��B���	���Ж���ꩇj�8M's?h1I&��&��V�8�(��>�:��s	x��x6�>�s�*C�i.Sa}K���5�"���4�u�޿z�]]�;q�(_�t�)`Ҕn�����˂������6��üw&[��<���!̌F��#f���%j�STYƅ���xn�FvϺ�k����p_(�e���0��]0���[)����h��/���E�K�g��7������Rg�l
p1�=��j�h��HX�ڞ�4ȄF7��!��u�c����Z��ũB���/븬�Ŧ��a�`b�Q�Z�#'A�1�0)�:�%������m��U*���n�>��Ѡ�]�6}�z$�Q�w�4V�y��{�Jy��iB]���F�X|G��łD��.��>e֌�М�Hҥ'P��V�MD�w�)�����QEO�o�4�[���^2��V�wy�O��Pб+Q�,���0��!"��i6Ӫ�yI�V�6w�f�]����,?z���bT���k�?)��"�a{�H�V.KR$����a �����T���j�FT�k�u���#޷ADP;��Lg��!� ���:�{�~�T�B|��1�o��yc���j]x��;�l�4�b<bJ�E��d�(��+����Qw�[i2��m�i�����Z�~�n�^