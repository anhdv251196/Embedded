XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������1aO゚A�L���|�Ҿ��K3u�_2�F�x������$��N����;�:�$��ll����_�8�U[	�Ct��� ��ww���K�����^�r��N���.�'����8��"8+�@�p�U�d�Òn�|��3��e�'��m�T;����T�! ��,*�fO�;
-}�����#	&3�^����Ǒ����r�=�I2�b��v#�[�L5�*�B�8p��}���1y�"Ԡ!�k���������!����Nyc�^;܇y����5���[M�޹�O��[�G�%~����[C,�D/�Z��#ǵ�V�X[b��yS2�&��"]L��J)"=D���w����g������X�Ý���9��	T��#K
��o4�|�+Q�˘1���g���e�\X)�(	�=�g��U'q��%t ,�U�-c��QO��z���S��'�\�9=� ��q�*��
_��G�ף(��b�i�4��_�э�����NB���x��\�5��B�S��e��[	��NܷV�NZ��Pܭ�Z�n���O�T��d���菱[��*9~�t>s����1�/)�ώx'�zZ��9��S�Ղ���cQ������Yv�}Q��T�q���̃�^�N#ov>wh��ao�Ab̋��� W!�{��B�|7E�uX���5s?4�^��c����d'�`v�>�6L3Dc� �?��Ƴ�f��J�3�xy�U���ܒ��XlxVHYEB    3c92     900 w�ZU/>���NѢλ�xt���� ��(h���\�,q���j�S���/��0m�l@�ir\�N4��%^:�̉9gǒL�O����)Z�	����;|Aإa��J�<fC���_+���l�����2V��A��>�.k)o�Ҳ�)�ڟ�b�:sGXzL�Q���`0[(�.�p�&Y�������[�H�'̌��>����q�F�� ����Wg#o0��F��0�U����U�H�����)T��"}?�����B��5U:HͶ˻`����d�^���p:d�O���wwAg�oX��h��nb��ͻED�i?��N$C�����W#n���}ⓓUk�<F0��o���3�:D��R� �u�b�B��n���̓;=x�.C�X���k�q�jOTsb�T �,��C�Λ��Op!�Ч����� l�{Ş�zQ>R��P]Nw��R#�]z$I�8b�f�Ø�a(DX^���w�,#�)̴ԿΆw��3�pac�C��E�mVt�ڱ,P3�_ŉ�����vyT�"��/{�2.{���*s��2"mg	����>~�z].[;ˠ�����	t�ͺ&>�蹸(XAH0E�Vg^�>��b�o���]�{Sz_\���م�ڠPY��97�25����m�2׷-���n �?إB,�5�|�����ɤ�ϑ:��^�c�hi���mX�7��s�>�$_,��8(��z�|甉f�͈v�]�r�������bΌL��Qy�H�l֜��Fm*8��9I�pn���t��P��ܿ�k}�Z��{���3��<U��,
0#�!��w�׊�?��>R�&�"�?E�R�	҉�]��};�t�!L��_�rf�0t�ڥ~.I���z���ד=}7�O��f]���B{OvĴ����� �7`�%���O��-N@��8�2�-�;��j�a��ˮ�ry=d�����{9�+ρP*�-6�OAUЍY�c�GZ)��S�C�ė�����nl���
�丆g���3�e�̈$�[�������J�_�6�P�i���ޝoIHt���]=W7х�\�'���r���|2��	�&�,U#Ԣ�ʤ�Z�S~Al��3>>�9u%�oٜ�9������0XT�ֈ��6,Z< �k�%ێ�_��w��*��]Gފy���#w�����9��������=72Z�Tyj�w��/UO�T�����Ƀ�V�
e�~[��0ɯ� ��R&�h�8[mq �wZ3�u�6�K�5N�O׻P��#w��!�1r��q��z^�J]�6�`�Ԅ�'��+��0����dY�̕R�%9��Ƴ�oos��%t�jrij��������A�a���딹��_�T���:.�!��S����a�2}�GSzKܐ��a�j=[;��z�i�ɷj���L3&<)eҺL2n��8����O��.��43b87�z���pz��t|h*T���#q��Z�Wה�G����0� Dʈ�e�?�q���W�|�5�8#�mk�J�X68'���\�f��!D4��$)��q�~C��e�)Է�+yպF����<W�c�JrK����bB<mO
d�<�/�c�h �`g[d�&�+dg-�sQnT���כ ���ogx�$v?D�E֚$��N�Ԑ�ʈ��/�
�n�n�������f��>���uu�%y]޳4�b�%�:4�c�v���C���Q1	���Ulhvs�[`s���<J��.��{	��+@d�L4z+��G,�	��H���MZC��ʻ���� ��`Wi�̯R�]%q(7f$`������f�Tj6��B|� 䇱�ㅇ�􌌁:R��F,��0zV�	���o*�B��X`��]4�U�V$�$�`�M����U�7�����Y5��A��Mq���S���ťAv]['���0	�����P�r�����?
Z�W,&|=�g�Kh������Tں���abJ���]!1�%Ɠ�n� p��͟"�4�`IiD1R9pp�x�8��<M���7���3�(��Mq�(���}"gS�H#k"�_�fexB=VPp����m(�u���<���˓S�_	|:�\3���bк���e_�):��*4��cYπ�uz���J��h�^~��UF-mM��+�Nv�}uk���XCF�����J�����ͧ,Ђ�����5�FZ�Pړ3�E�r�4]��q(�ZA�{�~~2�~n������n$�*�
&��n�I��>n�!�&.��H#iě8���c'E�~	