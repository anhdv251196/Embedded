XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��~8�n��Yd�T�����z:�o֭�䖤�9m�⽕�ϸ�t�'�Ο�����Ҧv}R�8K��X��~���+���)��/�a���e]�q��Ãp�X�_�J�������	/[�,��KHLH�b�jQ�Z�;�t��m�ߨ���m=)T22����RQ�n�*c�Yʸ=�E����ߢ(Y�k���� ϯS&c���s��$�خ�Z��6c��q���߾�Υ�ϱ�����q@��7Ä���>?��j��������y:����!�nL(6Kt��7U\�(� p��	ۚ��-|�D�,�P��<���g%��{źסBb�w҇b���<L�Jg"�y�'�v�����d�%xټ�H�"A��֕L0�ۀ�� pE�'4����_Y��[`�)��c��;Z���j��.�Ɯ�\T���#����`�Q�]��� �,�*�z��{e���U���
]E�e0c�YV�Q�E�$���n{�2l�np�V��aD��幠n�Ű�5t�����{l�T� ��J�`BO��̮f�l��7��/A�������4_�1.N��U����B�n�������(��։E5��vwc��̥��䈮���MZ>˟���SCfg"\�!ǣN���1�twv1��������ZPO�� nW4�b�q����n�0���̂YI�l�rA�J�o݈��*w��v��DZ�`��S ɯS�X�aK���1���H�D��L�Z�t�U�w�k��y+H{F��R;�)�XlxVHYEB    1047     4a0����������B��͓=,a����Z�4~��I6{E(���^���%���C�f���a��/��H[���rP��$a��2��@UdB��2}����;Y�f��Zl<2�X��U���@7� �g����Y��;,�}�{N��n�T������$���;6�zM�NHݢ�KI�g��L�C/�T~����	:����.��:n^��gԐI|Z
E�7Ю����h_�\�^���� ��dxӦd`fW�ms}B���T uwu���Zw�24~gSV���r>֯;I	���y0TQ\���].O�9č�\˽V'��>q���#N����<zf��C�#엺�,v`&x�ٝ�K�>x���Q�-2;��J�Q<�lA;Q�S���>�W�_~jv��Um!�D�'v��ڿ��%d����D*( ��Q����h���¸��3�$�O�n��gg�>#��NjO0K�'9��o�*��rk= �S,W}� �賍"d�6Ø#�KZ����9�oVNt�"�P	�����.���B�%115��F9��}��|%^�����N�?F܉�����vk���e���` ��Ю%�B��w
��^�=��K�&	~�"Ӹ����g��w��~T���\jn�[��s֮����0ê�[r"��M	���~��<p-�ێ���l�v9�"�C̛�����P�-A ����|hј2鈇���2RϷ��R�ӗ"!Q5W�>���;�� ;�1�����L11��y��|-+���47h�MJ�f^T���Ѩ�q��P���5u��� ��v�S��E����R��*���f�)��A{'/��x�T�L�M�$л�U���뽭������k����0'�
5Kf� K!��]�b�D��A�RL��pxK���K�ve`.ͩ?�Q2�e�~��|y`4C�{�<��X<�1�(|`�eXG��4����C�4K
�1�$(�<�z�
^4=MO$�BG�������a\��D���2>o�;	�Ķ�I�`#���e������8YJrJC(�C�<�36�NnC�I���*�����Y�:D0��r��>{jsq����(!+�UD��q���Ǒo�3B	�P��GB(�	�������I��`�2zh�]�4���^��yH8/�ۨ