XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��(�8XK_}�e�\�<�l���G�q�a�i�ͬ��[����)���h��i?�/�k�vX3:�E,C8Q�����;�zaL��ʑ9Z�RG�6-B��X@�c��Y}ܮ�5�!��� �ߠ}��ρf�Ѽ%>+w��=S��vz$.�#����>�X�8)X��H�9ӗ�w޾��%Ff��8s��8��7!�]�) �e�ER�1��T����2��	D��5�!s��
����_m*��ЬqAM6/Fp&��[������:��o�M��iZ��l>*����rD��������7���H���l����9@J�<t�]X�M2�ҵU���u���/�u�D&�1W���o�F9M\��.<�e�:?�l�K����a	�?gB��Xj�Զܢgu(�z�!a����5�{ )�^t�Sj�^�^���M(��,�e�7U���q�`�,�0z��հ-4�_?�L��7�k����"|~�|��7����B����d�N���_}	�����L�ߊ�1k�g8cπ^LQ��ݮS��%��(E����oK
�����Y��r��3�������\�x���+�;wO��h�c�+�*۔d��/�5�ZS	Ml82�dm��!,KQ�𒸏IoYm�r--���hc��kd��d�!a��]U�'{�+p��m����������΢�:�:+��cBg��{�w;zU(�ѝ���������<̓�.]�����x�;9�&�Pu�t���Q�I#��or�IXlxVHYEB     730     2e06>�>"̦��I�B���y��K�B�Ma��(1%��ғ�(r!��^'����ɤ�|�I!)=V���p�kE9G*}�f
�aմ�y�z�rp#^x�\��u$:��aw�fH�]�w�6��W��"N�lY	�s.ЯߠaԴ�E��tu���0�i��6.��@=n.a�z�nݤ�Ϯ2^��d �Y-L%  �z�����}_����~F=E�x[)\T��A֠�b�w�������M��r+�c|1��axARx��H���A��'G&|�g�]�X��r&�x���h����_#��X�'�K2����^.H��$��|���+�CdkJh^�!�a������&���ܙ�Q%�B!/XTR�3�\W &�([obG��ܲ�g��x����K�a��@�P�-�p�<��`Iȋd
j�ekaײK5J���5C���"�~����z�/�}�G֡�"��Yz�ʱ��� L�BGV�4S8ձ�s;��fsuqy���|�5�,�n*!U�(�E����]+�������ڥD�/��3��@�>�}s`�ڛcY��E��7$�k5g�ᤠ��c��/����cb��"���6�O2V~���b���)�!⽝�ʯޠ NqfYع�����2�;�
�'��ֳ������Ȑ��)ރ���۪�^���^��IN�nG��H��M(�y�:B����������%!�