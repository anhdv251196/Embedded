XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��"$� �B|� �{���9���/3��)"�ݏe�&�� [�)�ڥZXbZ�7���~�)s97�a������_�t�Uլ��	t�����%da7� %�SS�0w�f*��I-�Xh�i��ׯ�䁅G�3�<��sa�_pƫ�3��� ?����6T�D��m1pX��arx��q�q�Ξ��AOlm��)�/JL�>�l��7�:9� �M��~]���:�^�T�(��T2�ZΨ(��k�X��ɜ�^��!�'u����-��8����	��ػtSP]R�sj!�]C��C�޼���[VyZ�[	�O�۷z�!��q��`��D.�"��έS��	�l����
qh6EkQ�`Wj�Z���]��K��m�HUqv �+Ā���{�׬I��k-VV�C_\�a�|ޤU�ɂ�����,��t12��Ϗ
�#���8�^6�9���c��2٭�FU�9��/��P��${���;�:nF8W��0�!#�8g�(t9I��*��ᷥ@�j`B������]�ɖ�L3޳[�ff_{M����ᝋ�D��aѭ��Q��x���@g��N�ا�8%�!w����2�;K���	Tse��.�Ih�~���ΏO�����^�xwφ���*�a�$� ��-�;��#�Lg��r ��l�����ʡ�ȅRWf��R=ܛ���g]=�I�uˉ�� ])�5�+�x���5��נϯ�V?(���$���U��P�9�ח�qn �Ef��/�sզ��< �]�XlxVHYEB    152e     580�����Dϙ.6��6s�T�zO��[���jt&C:�Gޭ�1���a�Q!i�N�ƠdTs�\��
N��s��ֹ��� 4F��W4��HWE�r�8<�ϒg|����&P����Y�|���-��o������p�)/`��(�x3���l:T.}je��C8d#\�d��b��X���q�l�=v�1m�3[JXv�޼U���δƘƃZ��0��Z�ޤg!�̚Ce��Z&͇a��4}�L0iS�2c��>?`��tUN��ͮ���
.����|$
G\���"�P���la���M���`
��y������%s�bɿ2����p�lIS�'9�-�����{5��?�bl���Bk��R�;/�Eg]��=\�XB�-9�⢾@�W/���]�Qp�	q���lAf鄾�����v���Mņܒ���͊�O�����;D�k���2m���.�$�!C��I�od�1?S,[��`����˛?���l�|R�>B׭��7)�6��濑-���I|xw�M�4C�p��uE&ݡ`O����[��̐��W�c��ƷE��ދa7(��mQ�����`��ml�>��A��Tb���ɘk�1�a�p�0�U��S5����Ա�Y�Z��ǽ�XwGP�r�⭐����rm���4bd`���S|����v�\���Lѐ|�+٭���|{~98��H�<�� �÷����h���������暜��������{coiI���k���>4���'���>�h�a̻č�_�i���w,�-�K�3�v�E4BH4F��.�>�=u�{t�r>�`%Ҧ@��=��F�FȜi�8��rs�+�^��}:�ǻ&�R����'��?��FD�Pi�����N���2Y!�\�� �4��ȝ�"�{�4~�d[EH:0�K� ]]$>
�-ԋ�~��.�F�q(��_�Pp`��]�r�砅��S_K��q�}i��IƟ��L��p�N�$D�H������6�V�K8�;g�dn$��ߗߊ�d�	P�}��0qn��.��[����c좘\o�q5���l6�ߙ�J�aDT1u��dĂ�B��5��2���Y/
h5(�"w�E1n�B;�z�+5�g\�c�J���?� '����#�8��X�#w�i��uu��Ͳm.�-
*SQ�N��c�5`ұ��1�o�}e}�|v�`���Wr���cCTbG��Qh�)�:��>�����aZ���6�L5r.�e6˧���ء4"ʸ�~�0��b�j���-�#�5m��ɬY  l�:�(}��ųd.y.�4ԲW�=@�5Bt���u�˞B���G�-%�I�<ѭ��{x��B�N��y&��t������Y�8������8NR���