XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����8�~��W���ddY��M��@�6h������ڠn^Tz�hHps�icя�L�8u�'.>ܤW$�H�6׻�y	=�����1�>�3P樏���6P]&~��ސ�g'�ڒ�;��0�!	�i#av�&$J��/���w�f������iv7��%`Q�(��2�c���5+98U�<=� _L��~���c��/�2��g�����d�^�x�)�B)�����1������6���뗕���t�0�PO�����^�͐�#��%��GMb[����Ha��)���nz��D��qEM`1_�N$�F��-��m0�Rw�+��lJ;�̸�]=s�=gҋ��h5J��NO܃駥�Q�|�RY�]O�͟��'I�U��E��؛{�|nf��K����0Ӂ�K&b��ċ�
��Ɖ4+��υ��"5������T�0i28��,��W�����j- ���QE	J\(Zr�iί�ݏ��mEW`a#��l�C��{y�t��?����&������d\]w�d�X���X����|ð�C�;���aL�*�Ko�g	�*^�dcC�@�Q�L�Ez�2�Dn4M��r��'p���e������rĄi�1k���H�&P����f2�6������x��������;r�Pf���|,��k�<���u�UN��s��
��iaJ��P� ���4�,�;��I�XD�����C��v��?Վ$}!7������W��\��G�-�eXlxVHYEB     a4b     370�%��'/�)(�;��2y(����!ȒQ6u��o	
˖�d�<��3�e���A�bå�p(K_�U�a(dV������@�
���)�7ޒ�pB��cN}� |<�쿓�u���98%�#*�WkX��G�35x�W���SW��H6M��3<	Da�!��-Q��]�;���h\���K�e蓀�f#	Qӧ��5C@j?p]���8�.�;G�{.�Z	�G��B�:�����C����;���R_�f8_�W�6���:������y����Is�_�<e�}b*��5l�����?|�L�Dh-NЛ�:�8=)=�O�i�63��������f���~�g��	(*�Y;vu)ͪ!c����Elӱ����G���Ww]�)�g���t�'�'����e�&QJk�zS���v�[��HIܜ�����kI�<��hb�e'�u�[d<%Ba���+��eהpb�$���zitQ� M�+Z�\q&�:*K.�����N-S
Ҙ�Q�P{�
) ����(w�@~*����T�E�I0Ϸ�_��(��	� K}dK"0���t��{�@��x��"TVh�yȌ�eqR�����}�N}��Z�Dr�d��́�:&@�H��M��b�FΟ�렑g�E��CA���P��v��q��YЕ��LS���}�O�L�6����w�O�9�����P���^k>�}���F
�ddS�#VIrR��~ ���8��,	ۯ��a��'3� o������~�gށ@M�[���muUA/IH-�.���>�h ��i/�yW;l`�2!��;�\4\�=T�\�:%�&��r��$A�Mi�<}f��o���@5�x