XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���b�ۗ_�F0��j��i'5ε����Ň'K�t������RM�S8�vU�5�6G)= ��(!��b#���/5"p8�5	�>R�&\���ӧ=�G=�!�z�_�C��*^�k����ln��%��^���n��[U�"�a��bt�Ib��kaOW��<wO��C
��s@,�Q4���0�2�"��a�zF��vCL�BLF�E`�6�`I���Q�(a��.��ؓߎ�eD�VC���Я�Q����W��ˢo/8���(�&���F}G��p��x���Z�(Y�ڴr�8�L�[+1�3����S��"$҇!��6���?���K��2��nAB��~�|�*��~��U�9:�*��Ę���������Cv3�����Q�Kʖ����J߈�K4�i�x�����5�8=�����dM�k�Ƣ�q�~�� �����͎e��!���� (Q���s���2�x�G1s��;2�i�ӳ��3�-����*8>"9�nrO[TN��PN�#E���f�ݪ�_H���)o�l�_�ÞW��3{ߗ�J�P.	�U�y~��3��B��ͥ*}���I�����P�����r-�q�7B0H4�̑�C݃���r������bא	j���qx�U@Q3	'VV7D��R�A�K~�Zn)�aݸ��Q��g�%�	�/���)窿�]N���2��J�b�A��ϖy卤�Nd�z���r�e)�'�;���Χ�j�6���u.��qpC C��XlxVHYEB    6fd8     c30��@L3{�
��m�_��(�����i�'����IY
��F�����4TY�T_�d9�Hqѳ{� ��J�ސ�@�=�#Ty�?
���K�c�=���G���=̀w+�>S�%��7� g[(�	"�/���#Z���5Pk��d*���&#� |ґ�M�9�Y�p�������mF��V}
�Β�B���ݧ��a>W��dD x��{w�� i�5����s	�J�-f�u�r[�m��"+�Y�ׯäB�~rOt���+�Q���\�q�Tz�� -���-���� �dI����O�w��.�x����H8|.Մf�@A��y�Hۿ�K�Ҿ"�C!N�?`�Z;�F��N�a�L.=D��{z[�,n��:hU�/�YG3n����s��22�p7yq���Cr��a
)�3Jqx��xxn�;8��n�#��\Qy�T�����l�g]˶hZ�&�6wz�FG�%�I5;/�#_�R���[�-ث���4Ȅ�$�'�NHgZ� %I�~	�v~��c�hDrܧ�j���Ci%���LA��!�9���j^Ħ%��2���N���(��Qx/�W�|M�Ѝ�;˪�ge+�ȓ�D>\�"�/og<M��n�Գ�5I�7�Kx	H���xe?����n>�T�Þ�c����Wr������t�iV�E��-��k7n��x������횕��\�e���n�zl�e187��1p:x����¤��	J��ɾ%~��V�'���ޯsN|LLC[���4r�~D��7'�?��$%K=mG�[��8S�F,JX��ed�q]��?��'�#`�p�Lf���s��Όa'K�X�L̅�_N�)�B�M^ɲ��i�j'HFV-�V�����;~�_݅t���7ʡ��/	�e��v��)?tC�(��j�gC�6�[�jF��;ݡ�V02���yj�0��Z�br:�%;��Vx�>u����
}���{�d}(��E�t�/5]E�`�5V�q-A:3���j�Y
|���;������߈�=�Q����ݛS�=Zuq��aR?t� `G~`!	f��s�0��%�K&C �Y�����>��~�y��7*������ ��-�;�3<��Kڥ��+�w�y�r�c���P���C�@����P
x'�v���J���~H�`>"2>G~5i�EH�D�tY��gћF�O�ةt��O�q1 �[b�k�h��3� ?ڌ/�m*�}ov��`}�&�D�`jB��k/�@V��E�$̬�P��O�Z�?\��nt]y�p`����p�N����$sŘ~�'Δ�7ZhC0p�����h6 Ē���]w�]���<�Oe���3\t(��8C��q����!f�)� ]xXޒi�C��fȽ$c����Vۻ�_�B:t� ����W#Y�T�L�&��Q���XGfO<fH�)<J��lFgtWQ䞖c ,��cx���u\�$���M��v.����\���T��� �_�d�L0e;�a�1Uk��By�S	�.OW9Lby�O�C����F�7�]���0��"=�>Ftl�c�?8�A$5L��d�0�бF-�������e;Xk<I���e�ͷ",ZB~e�I���ePvC)�:l�dnP�+Q���3
��"'�����Ѐ)_�fݶ�1R�zȘ�q��)f�U��%�KIiN_=�qO����C�Tq [2Hs�:��͐⨮-W)�#y��d��wW:enz������ cLC�AG�mWw�t�rY¦0��d�rQ��]nQ�x����Z��ƶ��z���ҧ����j��;{:o�\E�pn���6.�|UM��&�ڛi!�|XVp%����{�i�w��f��Lq���#��	9]ޗg?w���rV��?Y�h�>�Hu3q�:[��e���joE�v�+��{�`ĝą> |���tt���jp��T�Cb8(�;��|�&7�$o���w�6۫R�#������u���Wl(��<�PP��K���3��Ś� h�.x�`�yh8�)4�A���6��r�h;�����Dj0�U�/�(z��Z�H�.l,��L�%w�LC� 6xUvv�~�}1��푱��J{�'��2�clBf%��r�Y�d֧�9�����&���[c���Ӌ�����ER_Z@���Pq����{A"	�f\���_�"�^�p��t����ZI�k��F��o��7O�B��gU��M�=�!���YVxʗ1��� �����P.�$�B���Qܳ�g�mbo�?�E�&ޯ�+�p/S֭�su�T��&�K��hi�M)�җO�"P��t;��)<�<S?q@M�z���ǹ���F%k��8r'C�&%0�����	o���vG;G�J���uC�4@�`�j������I����K��uk�Զ���/�<i<"�|��[P�%��"��0�U�@���:H>������(�I2�j���{�h�1D�Y�^�!�IH܌qa+#�BKH�<k�4w�_�5̾[	b�#כƸ�ۅy&�P�_w��^��;��E=*�#/�C���a.G�<�e��q�n�5cp���4%�}���@��]�hxW�D�-uˌ��,��`0�\'t[_��{4_{��&�֥�q(�^}��٠��0�X`{Az�J�Z��M��>}�g���)�B����<ȹ���!� ����5�4�Ugp/��QFt����h�B�`
m�<���an��s5DnMfw������Us嗤���@{�@�_�!:gΥ����GyT�_A�q�4���!�衁�o0=Q#��}!��AW�V�t�07�Xs^����ݥG�;���\�egdˀ؅_C���"jK���/׮�6A�O����B\�}�,����+i��f:�u?�<��dW��ԧI�;jw��~t�v�R�p��!ʘӀ�*g�� �A��k#��i�rȻ.�j�6gĔ�[�p�Ǹ.:~ �%��u��P�i��u��y���S4/�Uq�����D��hU�	�$T��QƵ��_C"��=�v:yq��g�ʌc:�[v����<���	"(�K�h��:x�!-��j�YP�+��_�K�