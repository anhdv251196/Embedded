XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����j�Ӆ~.r�Ux��ӽhB=��G���ʚ����ʄF�9�O��Ʀ�%���cs��U�q(fk��2W�0_e�Ԙ��%�p��?���N�z�A���Ko
�ǦY	�]���nFEԃ!�/|GP�;cǿV��������� ��oD����h����t�֢ᮂ��K�I��,ְ�\��d>i����V5�H�{���Ȕ��g�~�Nܓ~�v�4A��mG�??D�
�;r\�W�tC�=���������3&2e�ܠ��B����%����Kp����ψ���:al����6�vTx���Y0�F�:閱wjDFL���8�]�����������7��NP�.rd����M�z�������^���3�L�;1��\�ϲ?�Y*�hB�o�A�B�(39VJ� ]��X��G:�D�<OO�sSr|@�z�Ӭ��.��%��"�O$�@ �V���ݒY��>F��QSm��z�g�a�)�2U�\���s�^,���,g��+{�vc�	}�	�.f�A��0��Hk��<�ECO�M��-��t�IzDvn �n�]+�d\��m�*O�#��=
���A��	>�
�"��:"�G�wP��:��R�J`k:rx7{��BZ�ٺа����ƃݯZ��%�Y<A��п�2��	
��:HȚx)����I���@>�׼�P���B�Uh[\M���"�e&)���8����W ��dd@�H�_�*�ϞB&��O���@XlxVHYEB    6d0a     be0��i����	���.Iq�#w`,�4MV
#���x2Y�!�K�%���nx�Ш�)�ե��j�S��N�"�<�׃�<��ү>`��d+_��b�.�=��ϲ��O�4���K�H�N�����FlW�
�L��0_�1ש���32�EX���c&t$��q�`�򽕭q
o��N�pШ0��VJ����}.���p|�)/ok���
���I �:H{dĳ-Q#8�*]<�u��x��mN�`��=�
�B�z��9��
�¦;�$o�}�sR�4}� ��C���ۯe�MX��q��s����:�,�r�۲y�w�����cɢ+��h�>�|��:��R����B�1� �,�N"������eҭ?Z����OI���&~ًs��NB�L�qHC� �F�p�K3���� �\?z~�q��/(2�\*	ԄoW����WT���L�yJ�O>&\�(���0��h�ݭ`{=��C٘Q����̡����
�����@��|nQ�2D����f�DKPl�q���Ƶ��%A��F`��QB�@M�n��aY��'2���<RS�_!��pFV�D/����&�������P�v�K�d����_!��[�1-�-�M&�v֖`��z��h'��"�h
�Q�W�"NW�T���m\S��i�rC��������@�v���w�jU(`�6a�0�����n�B��{��h��3��6���_��5@�@�I��F�Y	|�bX� ����"����':V�����J�Q��"D5���zӉ�z��?���_CUv^�iH��Kr�m��x��U] �R�E�2T�<������w�+6��lȵ�]5:��1-A����b�ԅ�����_�Q�*_�dm�o!��m�`6	�#�G��ȿ�.����͏h
]c�;�W"�P="U�����.k���?V���0��wq	�'���Dp)��|���Ө�����;ֵ�`O;
��'�w��������;z�)p��(��_�GfG-�zM�%����}� D4�������q���cn��Hh��
��b�����N�G8�ý���x��r�t�����hY��]�)����K�tO%+�S�N���.��� �
�%���+n&�������������f�.���y��t�w�Fee�����u��Ѓ��S^��lo�y�t�c(��x�y���Ӕ�P�_�.��z��3W������f��iE���=U��%RT�vQ�8�����K})��r�؁Z�_�o�&F��]B����|i����O���.�i�cX��U��y^�x ս�����h`J4AN��b+���9v>���L�㭗��ђZ:�SM��d;�NO����gRF�ܑh�� G2v�����Gx��B£� P�!���r���b����~3|<���BO/�V�4v���>;�E�{(��=�s�݅�{�R��tI�6�Ƅ8�W>Szppfx�=��q�HJ���y_ ٠9|���n�Z��$q�U(m��%m �żS6�C���_c��f�~{�P�̈́�
�?��	�y��4(�<��V"��e\�AS�q5È�]'����� ��EmoOu�a��o�$�د��ڋA�;��W�N���� �\��Y�H�^����$����O���(�����^�?��W�K��䞣����}S�O���'�t~u��{8D��	[N|QΫ8N�5��KR��!��������Z�&��	!�ncg���~�� �&б3)�:���C$ǧ�y�u�Y�T(S������B/�,[��~�Dy(���s�"�5�����,���;&0�X֪�sfN+d/[�T�6n�%�w�l9��]o=k[F$o�_�,����1bU��L�{ύ6@����™-+ڢs&�%�ua�KO�&gGA9@���M���?,H~t?�E���bV[��h����j�h��qi�ʹf������rsFq�+�+W)�f�8����4iơ�j�7s�/�-@�ݗ'��kH�-</9�G�m���);���@�}v��A�[�<q����H	��J�#$^m*�p3������3���|���w�@��bh�=]�Ч!f&8A�qU:m���\ x�������h�����l�F ��n�A���I�Өj��DO-ѿ��;�4�bp��O����8y�'�L*N��{l�U@�$,��/�KA)ǌ��p%�=-C	kQ4l��FdX~���xg@�qD�G��Ld���`����I����S��1R��f��xQ4��_fbi�zs&�������78��ԧ�d`n,�?s�x糈kYJ80>���R�a�#{�]::?1�%�b��g0����$o~�[p��Õ�ۥBr6H� �+<�T�*�T��`GU��r�Q�fxnRj��z��&r{W<yM	�S@�5r�K�G�R^��zC@.���/����3h������FN�L�����q���������d�����`���O�'�"���T�>61�-���,�ٻ�؜��C[̻Rf��_ =L��� �r3�z�%U��s*W���צ�T��ݜ�x ]hwa�BQ�gtS�~�O/6������L����&"�{qUlM���
����ũG�L�C�&��b�i
..��`��^�ǟ�?��S[*��"�,�9T�v�,�+xG�*d�Jo���o�]�j¸��׼�^˹�Y����Д��OC��ŷ|0F
C�J<.Q��*� 65HFS+H-$�/��DyN�a\������9(��^�*�$ �s���Sgb���
�j�0�y�7]�'�e,Mil\�d~,���d����?��7�(�C����~j��͗R��-�`VUȆ	�:0��{^��%� [�X#6B0���$͇���'�F˅`�l谫ƙ�!Ծ\���g�w��~��	d�0�_�<,�\�Era�$Z��.쎖��}[��0�ח�g��������0�?h��.%k�qk�!���t