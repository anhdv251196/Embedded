XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������^o�RȚ��k�o}P:R���D���[�6xy�cM�25����:���Տ���i�aq�����'U��&|���;��&�"_��~r�baY���@���A�)�`���as�-��;�������g<��o\����RM����&Q�ߤ7�R�-6U���T\���Ŷ2��\Т�B�K��sRv�-�á�6��S� ]Hۨ]ȼ����нe��m�%���M��e�1
HU8�GF-�w8[cVp�Bb�=���;G�����p��ʹ7�W�	B��e%
e��'���h1Ӄ��X��P�q����x��v�~�g �������Ǧ�-���׭tj ����+�ST�^j@Fa���L�������|m�3c�>��٬'��C�^,.���<�ܚq�ǎ(�F�~ g;-�T I`CזN��$1r#h]e���{&8�_�Ir�p�&�ENi@��<	�O��M8�#psUr�����za�!u5oI�Ip�Y�oYI���=e��X6��ޫFT|,�G*�p�e���մ.e"�6��=9���8FΓzB~��l-�_iH}k�Uc}υC��_T0��H3�`5��ևq�C�$:9�e���W� v��e�`=�C$3,/�3���7��:�[�R�fFX�U��7�^�&Ht��pU¥�C肜h�.��p���1�b����J;}�}��So�ۖE��w��!��˵�� ���R�ة�lg�H�sޙE�t��j]���7rUO���-ey�t��h~�qn�S�XlxVHYEB    b892    1b20���0�6 ��/9�$�}B�1���WN��ۏff��/'���}R(g ��k5�#���x����� <H�dG�/��2��Ҕ7���o��b߳��g�h��1E�?aCJ��,ocL��&�#�g�o'� �'#0uC���w��K{��ĝB�!8�L��lF|F[î���p�qiV��!\�eN�R����pY��޻�������̔��"xCh�]W�c\ö�5 ���Ԅ	��0(��9������� �Q��e� ��+�%��k!��1�V���[;�7�Ԏ����������v)�,���O\�H��y�zJ����Ki��T��%��C�k�#�Dk$�h>�W�ä�֫`���?��?:`����������~�A�
4.p�����\�����s2)���{>� +j���H�MIc��wܾ��g�t�`��c��Ch�b�R�����A���&����P���a�ぃf��p���Z׭SS5�_����o��M�M����AH�q2�ˮ�4ۨ����6xJ*���>� �lez��k�&:+s�#~v�'���\ɮ+�eS����7vl쨚3��r�A�V#�y
\��q�C���YC�d��\�v�����W"}�-7���H�.��P�8C����8���繛|	R�;����~����Y2�Q��� ���mw-L[�as��Gl7rh��t��y,v�Tf'��;����Z�D��/پjy�F-ݲ7X�d�Êk�k�z
M:J�q�%��R @�.��������
�Mъ��N�Q�ǣk@%:�3U�pE�θ���E���6�L!h�9%@��ex��߶��}yڬX��R��E�d�u�6B���
�m�M�ߝ���8�m���_,>��#HD�8���������&��H=��֗s�bx��vU�«��.|�_Ύ�ǲl�j_Z\����OD�����s
�f��#��	>���
S�pp�G������f�����._B-�Uw\t��'�OUq-|�mЁv��;�xI[�<U'��̸zO���XC1ͫ׉�����mv��i[����@5F6C��^p������4�=�`eOK����e�y*2�Щ�$"j2�*+��Ɖ��� LM�|O��^�Q�$�:bmp�-�x���Ҝ�`1 S�_h�ا��#�$�J<a������M�|,����'^�<A㐚ϣei3�BU�����bb0�^ʁ"��E������M��%+��޼o�t`:�n�6���_c��ꠗ�ם��歒�^Fa��k���<v���/�ۑs@�=d캿��Ǘij��ts�4�Z"�m�=�'�Wک����R���M�4���.�+��[���Q�㝫�;��/;q��| d��v`Q؊J	�����H���2ad�6�1L.br1��0E��lUf�.^<�x?|&4�`v.��>�Y3OTo�^!p?���&^�m��:�%=d!�	?�%�������
ɶ�ݏC��l�H,�SLi"R���r;蹣> �$őzx[��[����,��+�T?�&j��/9��r�bH|z~�Kw������$�����{Lm�ڇ�v<eF��:�����;[^E�������e�0"�i����s��E���@�����J�����HИ5 �6��-��A��b�b�#J���9{�@0�y���2����R�j(<J\?�}����Ga"�xȞ{�;$n�*�^#�� {F����K[�s;o��/D�{"$7ܔ����jڻ�5E6c�1vM���&*�s1�R�JJZ}�K+ڷ�U����g�?=�qڮ�"�GdM|�I_��~ -v��}��U�	Ve�]��̈#����:R�q	dD3���I��n�<�/�0w���@Bb�Oh��8�'(��:�C�q�z��c KI����Im�r�C�}����2�WƖ���M� �Mx�R?��5�[�]7Ω^��V���i�=̿2;[ T4m�s1\�嘣��J��M4��+����`<ہ�I�"-׬�ϗŹ���.���%w&Bi \le#�k�Z^�
�Of�Q�4oU,e�{;.$��+WZ��pZ�~�PZ�đ�F�aTj齟�5�v��vMTY	��U��Ӑ4��y,��tb�W�#;0rH��M�>�����#ϗ�'y��5�H�T��9Mf�[�������g���Ј�#� ��7c�M�����{?='G���t�2�=񏔷a��Ax��d��J���4ꍽ�ì/cGGZ�SL���h|��z��E�R� I��@�+M_����1�=
?,�ت��I����j����<wut���D��;)y����.2\�}F�	�}3�p�(c��$%ӛX�l�<����se�a��㾾{G,i���\���/?}�ԛ����BǓ~Ё_K�=��b;�zr��=�ۈ\rJ�|�>�%κ`����=h��xo��IoC(�:&�%�Nw��f��T�bh��f��:��f�̈́%�E�K�c%k��-䢢u۠�]����?�Q����[}y=e+ �sy���dh��NQ�/��Q���^�~(K���.!O[���	��v���e+x��#�@�1L���9��)�qO+I#����n�K� eo����ʄ{"}��f�^����C��},���H9�������J���S�݄�K�Fs���.�N��"B��LUa�O�O�׉�0�0�~�G���)�6I��B�g�ۊ�������e�\4��gieq��e
<�hNs�g}���(��\�����;��w��Jz�13�<����=W	#�h"���R�A�a�E�a��	��U��� P�#ě�s/׾>�fK�pMX_K�XjVkK�����yc�xvN^��w�eg���L���%e�IQO6���E��WԤ��q�cB���<҄��E�t%K3 �o ���,�	خ�u�"<I9(�1ģ�p�Q\I��L*M2��+�^�����L4�!�!�M.ܗV�_K4!}Ƌ�8/�9���:�	��y�Bӑ��~��I@��2��b"�h� e;�<D�!�) ��O� ��n�쪄|YЪzR(['dA n��K[��D��x�C##��9�����E�V����>{G���Kϱ��|s�\<����wx�@�E��}L>��qʰ��,��,g�`���rm�¨�2��i���܃g�*/NM*X�Οy�\8���(�gD�X��7�U����\p�^��y,�T.�X?���bm��p��Ѭ�z}��RG�$���l�O@ݥx���'j@���Z�9�D���U��\۵�?���5_�1W��߫D����Y���u�J34�<���UH��*��i�'��7�%�U٨�;y���v���+��hRBPi�%��
�u�����>�±lĝ�+����2*�H� q�_y���w�'�D%ӥ��U�5�X���j�.�M����A�W�Y�I��X� >�^N�J+� I�<��xX��3���Yd�3H�'k���I �%�\1 �}�qȦ^������Ժ�@O6�yl��ͮ߿n'����4�lȸ�ՋNT_O�ar�b�q��7�ֈ�]��%�}UA<�KV���[c�9���S�(N���TƔ<d\�.��h(àg3(�Ǫ�A��䆖�cb�_�!� ۾�Z���&�w��p�A�+}�δuvg?��T�v�$@�6
�z��� aN,�>͆�����N}N���wb;�/1����&M�N_�L�CG��q"�(r���������.�,FQ58CF�W6�n�2d��x6i!�0��aV�[~��n�+���@N(۝oJeI�:��i4~�������я�������e�?��\�]���K�x��	��Fq�R�U����ҭ�I�O�&��\^@�HL�%�Q���xmY�69�0�Ɠ�Jo-�y����m�r���=)�&;q�r��W��.߅�"43���"m=��RY��?VM.u�kC���\�L��U_6�i�u;9o�,i�zH8y`���
ݘ�p7f�ڋ���a$GF�e��STni3#T
��G�p�����n��lmP���biY�vk�w�����d��F_K(��2l��7$�z�;?�=V����c�0S���&�$b�Ā2o��p�Zm����]��4����:�H��;�)��I���8��,��_��Mۮ�yS�U��VOfe�˝N�I��w`�zwװ�������j�����
|I�(a���RH��k�*����ԅbz���xPf50|�4v���2˅�6�;.먳rMh$�H��8���+�*)5X��mK����e��7^�t<��9V�.cz�A�����ئr�,h��8�.�7�	�C��@qd J#O��\C,�]F"���'$E�D��;wT�o�Y�`|���,�h����n6�}8����*�̟e�NL���1��ڡ�<���<�*wF���@(�G��f6�t���X���&ںv�'nU��|��42��M�O�2��2ȱXQ��F�7�}��z���hH$q�4!�}�������R�*�MyH�x���g:�~S���q���,q�j��A�����.��#K��3$0_�%:�g�{��"wsGK�]B�]x��h�]C@o]���"��h��Q�t���B���}��ۃ�6��f������i��LWbr�R�ow�p�D];��/�Z�����|&|:N�n���{���=�P����b<�H4.�C�Q��A���G- �_��6�D؀��֫#;s�:&D�TM@t��Vg�g#�f�	j�j�.y����Y<K�0���2f������L 
�Ț*��K��oE
ܨ�Ef�W�C?�'Ъ]ٳ�/���Ux����V'���Kb�dSX!�P��Z�p�W �7�P�,��:�m�y � ����N�M����6����G=At�d�.�U��p ��k���z�w��-�"�gG�):��}T+�� ]x˼�MیK݉l+�AG�����o�B��LLh�P���q���˖8�[��ҫv����c��߹w���{ѵ���a�X�Iv�@]��C@D�Q`E
�x�x��O`�i3�N��}�2����X�v����f~�+�	��r�Z�,�0 H�phs��H!`|+�xvr�0jq�R�Z���~%}ʃO���Ү�nvV������Q�p�Rw���-=�I��o�y�KL�"g�m�l�+1�.UbM�y��{*uLP6�x�m����q��н��D�n�qA�$'Ǣ1e]�Ĩ��s���(P�����%o?�TM��:����;%Y���m��pט�*�������p�[�u�+�^�7Wc��
�e�>S�4,�$|�x����\��O��ܺ줯35#Fޞ^�ĞH�?��b,m�����"�۫�Q�+��Z���S������L��Gk?R>pYd�BD��=Ńa��5�R��+�kh+�!w:;2A�ry �� �<%����}d�m6���Ҩ�����:��w��=��:�p����Xz��z������ԓ��/n��՚3�<��[6�1��i ���4�������w �+���F � )ϲ��X����P2���#�&(�Iгq��N>������f�fp�XX����E������#^7 �Xq�$)�=�=���$D��%@<�		�a]������>E:)�����*��pOX��z��$O.�o	��f���v�Cr�7'�D�Ѱ$R̤$b��o��;.�.�D��΁���Ɋ�ԃ�>)�.�L�������jFɥ��AW@ۯ2���$�K$M2V)��NP�߱���U&Ii�ѩR#.*kx3E��U|))�n�7��#����hBd����i�%�[O���� t$������b5Da�2�
���c��0�?�
=B����L�L �n�N�f4#[!%�|Q�ԟK6LA.���~8�+� gW��}��[6J<�������0��� ��� �d��g�to�Hz���1,X�a:V��$�BeI�}�Fٌ�1��?�m���ׅd�e�d���k*s�A<2�{f*�LU, �<�,�D(f�4��`r��od/�ȥ q	�z�?%�#�c��3�z�mU_����)&2Ki�j�wRL��TÞ�#�*��:M����ban�}�
�cB�������%��H	��6���EO9�Li$�;��˱����=0f��%7��?�0NN�+їóU���5�'e�?�V��!�`����#�e�u��4��pۣfi$�_�����
����j��¿�]<�z����%_��sj��髝�3.@�� �4~�+�K��c*�H�i 7��63Ҽ&�n�A|���h�~�I�+H)*�0c���ʆ�˅����pO��yy􃸜h�
13��oi͸�2��'�źa�<�$t���/$1�)q}S�,oA^���,z��%y#ސOyOD��)<u���s+?�Z?���oF���*t;V�˥K\x��seh�%�s�Ja�I&ڭ����b��UX�	��2��ܦ����s%��
�L:; ���x��9w���#�	������k��P��]�ņ*&4 �$��5�M`�����y��NjS�L�ͬ|�a��� �.������{Ɔ�_�r'0֋m�t5 3ԇ�{���6�[4�/��H�[�:ξ`�\�X�>QlM�mt��������z�>��QsY�u���$�6&HX�P��"}�9�I�x���a��`�s+�â��.�ОĹD_����u����x�,KB�T��L0".��J.R���u�k^)���ׯ�������g���.�	�cr��6�