XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����5P�.��*��_j	*�����^�^Y�%a$&ww�AFL���L=�����b��k�*:��Zz���{�6�8ٓ}�{쳌�/Og�v1Y��gwu�u�oR�G����������y%�r��[:�iv���-��<��/Τ���Ⱦ��k�&�T����2���	�q�&bNS��L@�0t����>��"F�iZ��N�$q��+���v�F��% ���f���Q�a�����ߩ$d����8:a�}�٣��o�}Q0K~[*4�M���9���
7�D�&����flu<*����	�[�3_:9��Y�������Ǟ4]4�p�n�M1R��맚��L�P���A;���&c���"s����+���Ħa���v���[��+��ʝ�1��h�@�ڡ�u��H<nOiD,}*��l�eb����X�J91����x���1Ɂ/�@#_��ݍ^��a���zx\�R�,�ta���3¿�TW��͉�R=)�x}?h�*���#��`X�n̶ͲCf��zF�^���O���f*���#S6�7��.��7�4�?���[�=Uڸ���q�_8��d.<vb��9�*�Y��VZ��E�0��=$�����A�%2	Nh3��wE���G�n�f3d���I1sA��$)lឈ�Ȉ�{� <^�|�W"h�֚X˻La!;Q*|�
����g���v>r��T���}Tp��	��3�"�=���o��*$�#S$�qXlxVHYEB    1046     4a0���(J�D�C�J�U⦶9f��\���0̋�n����]�����iVϫF�'y�Aty�ޙp��ti�J�Mp���63u)�?�6�]��TңAR#�-&�h�r�R]6��pN�p�����n�q <��d�k	<�(ƫ��/��15�ˇ8����R�j�G�k���i?���-i�M�2��3܂�Nx/.�Lu*�oʍؔ�y|p.���g��1�Z������oP�(d+C0e(����r�[?�,/��Q���AL�w{��؛��'%U�0�y�1]��*�ظ�������<�T⛖ ���A��#��P!��=7'y�8K�b��xT�t�(V"5�l�������n�c�Qrm�_ޞ1��t�i0�]��@"Sb�e%M���FcZGh�}^��z �;�0#�Z3¤�
�������d�����jB� �F��m�α>�%��DY���fx�:W	l�}�8E̤� ��l� -��9�Zw����Sju�4*zr>I�X�����2����B1��Ã�n�U�S2�$N^[Z@a�K����̡l�q�WQz���	uɼ��Uq�a݄�Dۓ} �l}we�N�����?q`�R�o��7�^�{��_�t����f(A+(���/�w�NS֤9�����&$������5s���������+)���h�;!��Fu���_!����=�<"!�젭���~m�r�??�ǪH��1Y��a�J{:��9=X�����n��e׾�����K�?� �3�~M��ab
�V�Ƹ�����y�(R0a�de����c��Y��?�a��=Y^ہ��-����q��!ßH��aU�����sw[wŧ�!9RXv���'���pG��`f�R�s|ȝ7䕳�3b�G�f��E}�ħTY�J�s����ec�EF�q���������G8���@���7��Z��p�J�yP���`�Ҡ=�<N�ֲr\���2=y�w�('6SUf=��|S=��(/���w�n�_�T�[�_��.������!D�����1�8��� 2���2y|���K뷯gLt_�I��\sQH��1����q�������'����%���p�i���-�Z�����|����߫oC;�&}���0���XQ