XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��R�l"!��m�@&��m�e�~����b�{��}Vf�����B����3W��W_�ui��l�h�C����D�u]Z�����v��XC��e���OnFz�(YǪ��+�+%WH��u��[�Q���rOf���R��g ��ˋ���Y`�=����,M-�t�J��B����tܝ���ƒb�$���� ѓ<"�n��au�'<��Z��R�*#��n,<B6S�0������=���?O~ѐZz��o�xU�c��7�WqN�
���SCZ܏�1�%��.�HN>��1P��J7��˗y��3*!��~�	�V�<?ƭ-��Rbч�r���+2�6�	�s�Rt�*i�����J�zݶ/�'�6J�R��@�e�^z[�<S�(s�j������};PN)�<N@Y{�������Y��7���9������R3&�Ǣ����uF��~�;�ռu����YԪ� �r��G����	
��J8�A:��cn/�����I���퉋G[[��c���3�UT�6��.s���G*��̈́�L���l_|��v���y�˻[���kd��<�#�H��=e4�Y����E��u�<�Y�Y�m.A�8����n�����g.z�eh3j�9�C�H�j����W�AL��(yc��@����7Y�P[k+����[͘�`f�#�h�Bu��Sk����n�9�y@l�
v�I�������,up�ѭ��VfhR�Y��������gXlxVHYEB     686     2f0�O�ް͵?2�Q��Ε��A��o:
��0�yk��@�@;t�=�D��&��W3e�����]jE0_l�e�b�rP�9Ъq-����'�y!�	��,�z�K=,u:J!��K˷2��$�8e4�MR�"C��?����3:,1�6+��e���R���01Yg����c��蟒1Y���mF{d
>�|�g�K�$�鹸6Rc����nCƣ1r�W����6��jo)��I�r�I���LNF�4���1?Z���vD˫�>��|D���ܷ�A@f�NDn���A��q���������VZ�<9(ĵ"��a�N>��n�}P�yn"����Or7��/���!��/I�����6��:��ڣ>�x0TA�u Y������� �C����Di�:�m�z���/t9p�u.���?��B⏿G�ګ��$���q�@�4+{�X�J�y�y�m�6�퐅��J����A�BZ%+������ʊ\�5ޏP�1J?&f��c�ݹeR���bB��m��,�t=�^�����C9,!���b$qW�L«EG�8 ����c~��|������9�ir�X�l{gm�L��j�΂�L�@���p�P߰��Ү�D�Q�I�=�Vе��#��4��4q�X�XSuD+�䭯Ih�(j��"7˧�v'�>�}�X>�t�	tx2��a˖����O<#��U���;&�̒�D�M��Q�NAE	�.n�Con��ɸ���!�T���p��