XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��B�b�u%�@E� �X%�s�z���.�7��	!�d��Fs\F��%c��d��n%���0B����`����8�[bil:�W�c��olO��������va�>��1zq3?K�f�t��pP���@{;n1��\��W�7y10PJ�%x�x��}��:͐��8,%�M�./��?٘�o���K��Zз"��l���S��^��Bcp��x��B��� Np%�v�V�2��S�(��d[�1�׵No��LX{�&"#z �.�}8���E�`T���D^^,���]�t\q�u�K&Xuיa�Fo�e���c�ͭ��.[u���͂AјE��~7��x��4���^��:�>ԏL"��p+OL���v���%}�(_�Q��ow�jȆ(��ֶ`$����2�K�������Ϟൻ����)T�BS���.�W"*x���>��	)�^q����pP/M�ȧ!0�'3 ��(e��貛a�_v]�h ��Q�{���X�s�����t������7d�AN�H����֩��S��E�Y�r*�P0���p���(+�u� G�(���nb�I���)b/~�;]�QA�i�L�ڟ|�=@��3O���nT�U�����2���a�X��ن��J�>S�R�9�Y[X�G��t$vg@�����۝����W�X
��_��_bɩ����A��}��ֿ-h���E���Ѻ~W���8O}?{�y��s��l���T$�6M;��@6�j�&Wu'r'��kXlxVHYEB    1d52     7b0FP�3M�H�	0��|P��r�1��C����\r�7�	ɤ�Ќ����E���^�RBߖ��[">e��������Z�4H0��U4�����Юq���M�u[�F��x�e�J�I�bAҺ��6�r���ǣ���r�aD�d
� n�W�Q�;��!|���BI�*�|�\Ђ�� =J�cO��'I��s�5.q�����b��V���M��Xm�j
A����v١��Șm����|���w�}�g^Մe��DH���2�B.7/V
W5N�sY��T���_=�ѵب�פּʌT��s����K��3OQN]AfPN��f����А����/Z\����
uI��3�5e��P�rQ�C�hH����ܜ^�%�s�����<"^˃,����G�%�0I��dv�ϟ���j��(�s!��9A P�%U1�*^/��D&��/��ЮZ_gJ��	�!�#��"�|��snԓu���]�+b�&�7B��Q�N�B�W.O�V���b,��;��G��4�GdF�]#�D%�/7�Y{���4�qR~�y��܃��%�<�_��E�cj3��_��>�*v�JL��c{ќ8�� ��ՙu}��IC��|����9$��rOY��is�D�&;�q�������t���p/��xu�XMT~T|!y���ۧ^��z[�r�B�W�Sqp�������cDL�]�L;Ls��UM=����{�ky�r��!�Vw_�vh�}�+;3���}��=*r��Rׯ�F�V1�lF�}�^�H�7��v�O�	^�o�/B�f���6
i���t�B|L�|S�t�^!�����i�K
�o�&��:�Ǎ�3��_��+ ي=��������_�X�9�I���cp��O���]y�Ϩ,���tҝ>�=4o��x.A��q�=w���B~V��9�>T��)�ߔ��<�٦�޺Y@Q��`ڼ��wi���M��]q۝�˄�D��<���$k-+�a�j�h���N�UE�l���.��:|VipF"��Ұn�K��n�܊�|d�Jp�1dv�D�LqC���]ۈ��Rj���^��T���F�G�H�ZЪsQLQs�o1��yT�q �mΎj��Ar�x��2�?���7NgC�n�H�<.�B����V�"b�,��a��t�w���w�A{�\��~�AJnɓt,�mt���������C�Z�0�\Y�8���M��v�'��%��BH^N��J�,Iu`�3�����n��S�`�/vq}a������P}ܟ� �<�b����F���W�-% klA����W��폂�
�ԯ0��H�(���R:�,�#�����Q�u[m��Y���U${����ðm�l��>�����r��J�\�D��SDO�~���<(�{��"9 �\�,1s�u&�K�(��ϰ ��~����S���L&儩�I��$�(��k8�R��
�m�@��*���iA���		oP!�9�K�^��\w���K�H� 4�`�.¶ZT�̟f��Lj*+t�"5T���)?��ih��A�hg}:�n���(�jQ?n��� �r��I�!Zx{�A�MV���ᛵ1\X�[#F@��l��ǴʜH��*(T��W�/�9�M��A(�c�m�r�ų�.�*�؀?J�&*O��t�����=PFt�tTzn3{�ǣ;���U.ܣ䊹�8��V�ʏs��ٟ����d�"�/��8H�hF���Ak�f�5���j��W��6�iX���|���Z���V����՚وg�Hl%��Fi��g.Z,��"�����Sr|M}��]�i������p��x�v׬�Xrs��@J��R�B]�C�<�][�&K���a������!ƬYt�˴Ƣ��@P���?�H�?��+C�φ+i����T�(�1��