XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����=�U�O͏��mg8P���|�D	R�3�I��R���/ڶL
ڥ ��i���6�"��6e+$�#F/�tٟ㦠P����ӯ�8b�I����n{<����	��J�?����*�s�c���S{����aa(\���'6 @-�6"ʹ#����B-$4�PI"[o�Ǖ�������pTJ�z^�d�+�|�����w!{����ǩf��P���p "��2��e\��%-����M��LN!��X�Y��-W ���a�ó�s�e0%�@�p��Pm��`|LcsM5v;`��$Ҡ��b����<��L��xɃ5�U�g �Y���rQ��{�3�i	W�vm��<G�%)�ԱM�̸&�/���P�Q���NЍN�}y�t�β�?)4��9�=X#���t�c|�;����m�} %"!�_.}���R��kz���(�,?.;��T�X]��y��)9r����C�;�i�1�5_���j'�w�G���N���k�(g�Ƈz���EL]j�;W�r�ޱ|B/I�N|_+W�l�RA�L���v���p,�}UI>��1�� ������x���KOVx{:Ty�0�.�\����cЏ���&�%]}�*1׃�<)�X�B�B��Y���P.��8��TY�x�xo�wO�׉��>�秅����xp	�擳����L��dg�-~�'�`2~���n8Z�?[P�n����r��^���SC���o�ƣ���P�c���&�XlxVHYEB    60e7     cd0����n�!�@�>e��F�$��_i�Cn��@�4lz�D��$�˵"kJ2�0D.°�t��Ɇ�����z���9؟N��f{ʝ�J��lN��ՙ� #��㽤 6 �E� ��pƺ�6:�Ì>�|�����Hp>�������@�Y�>~0 {ÕRT*�	�le�����"����m�/u�^�{����ܰ�,�u����K�aBA�����p���D76��t�5c����6�N<�n�2@��D�&��Ũ��kTQ���Y�۪��a#��K>t���Ґٷ'.��a�%��^�_8�7$�9�����ͮFW*��>�����nn�5��;#k(4`�5z��ڥw�hK�z���%F��}�Qf�ϒ[$.��ҥ�fި���d��-�X��Q�|#�܁Q�>z����1���I�'ə1��+Ҫ�P@�^�@�&A=HO���&Ο�&0Yv�-�m�BT�k�����%_yE�<=G�����!rݚ���	�I�5)�qfx�W��˰{�'&��z� 2�q�E�Ih�H�ϦP��m+��7�<·܁[j�F��,��a����v�c,�졄"�"���ۻ<(Gn��$����Ġr��rZ=�!�g�2�^�Z���iE�k�=����
��<�5"���G�>������ɱTc�S���(���~�HqA>�#�{���Oy���$et N�F��s%>�VŢ=��~0���8jӜ�c4��;7�h��Q��]�ЬmB`'�2�T�� 0��~zt�u��ܧ�˾G�7M�������Gc��Q�]�?�-�3�Q��BH�!J���'� �Cal�������ec�=8�	*���k���� G5�F-e��q\���0�Xsj�_F�ⴷI��^k�1�V�`@�b��G���(�ƺ(�3h^�6�01���~?:�	})��'�!J�Jo� 5�v��"H��$x߂Ƶa��?��0�6<]���D֩�T���M�§�3]a�9��
��4�+4Z�'�Q���"8fӉ�Fw��鵏q�b��%��'3E8,�6���s�y�C~�yPީ��e
��?��
յ��D_�HwJk5���`,(�p4Q~v@0�4����}�n ���	�x`]⤃X���������̺�n*u���YcU�� ��;I�'������4�^�"7#K�9{"Χq�6=�����рL�-�4��.���,��k����`5`��|X�ؑ>�Q�o+�xr.0���Z_@�� z�4��8 a�3Y�����F�nM���c�%�S�i*i
[��-�"2q̡����7��`�����
|����U:G/�{�߇�).��j�҈�`���m���0�%#k���Z6����,;����#�'��F_Ƈ-	��)�A"��v��֫��R!rʓ<Ţ߆��zH�Z/밃X>�^�{��7U�wʭt�G������×������r,���A[����։� 2��G_��N�W�U�T�d���	��f��T�HW�z����s�I��`�bE8]uu�����&y�Eê�ϯ���L���e��9r)��I���<7KćeG=s��j+ -iP���ޕƓe;�*裑��w2W`,N�Yհ���ajM���ф:P���4�s%�����'����/�i^�	f�ǌ�j�?�P�{B�X�t)l��sKT|tÛ�mT���ĉ�um� �x:}@��`��ݥL2��q�@�O�5X��WjޏT,�`iA�0n���4���r�}�.�����t�.��_,�+2.�ݬ���ւ�G�گ��O�i�};�2^C��m��@��q#	}j��W�
qӂ�61�n\��R��t�z�!N�9��K�g��Zd��6�n���X�S���6�� �jA��)�\p`	�������Q���$�ӭ�bf-�FUZi���ё�)�����Z��q��)*���Q��C+vl?�G�5��U��8�}��&�����޿�	�!e�)埯�g�������;oi�s�X�'�O-��}6����5�9nz��J}�zW
��}���b؊��,�ϐw��U�����R�w)|;��9V��6��sQ"��T4˲�a+,yr-���i�t�Ӄ�*�?��s�9O�0řV���&-:S�M/Bx⏂)p�e*�_d�R��ӧk�|y�S����L��N����V���E�l�*)�[�w?�Jk�ǑdN[p�̵��w��s՚����憒`������7[�Z��j.w"E	��O`���D$���M�ƌk.P8�F��@�M�k�G�"�1��%35�A}�#V[��bE�l�K��to�қŜHs6��_N���M��g^�t��k����J]U��#��Jj�-RU>��䔨=��L)�����V�;�eս�c���M��{?�1U>�e�iw�Z��G�~�l+1��L�2��/s�jr	+��")�b�8�b��x�?K��qfJ�;xg� ����2�i{�燜5�v�Ʉ��q��0�w��� Ń�c\�}�:�8m��}�GOr�y���۝�]�`�;T���񹳎,���w�]|�Q�G�Z�>"�����q�CW�����K�ZXP]��pj]Q-o1��&�th�
���]�^���8�5��!��[
�G� ������/�sؘ��NCA��Gaw<�7Ơ{4��b-!�V؉�I�gƌs���y���.��21��]d0R���(B�$�x
��_ʒ�co��3�!�j�
��ktoB�>j���^�E��Ƈ4gѴ��M��N��F�-��k����`���"��3LV�����Ĉ�ivP�zp���O���2� ,�p�F2�'�8�.��:M+!uC(3��L��lt���_���Є��q/�J?��4�?ēQ��K�����ԟ�M�����<���/}�>V%����馑w`�"`���Ҋ�_�����|n,�Ay��Ps;�b���N�S�1X��_d���ڦ�2)�V'|�����.`����	�!���y����������'�(f�p�B�5�ն�X�ٷ(G�*/n������,^�Bő!"�t�e8�2�K�b���N4�|C�-���f�f�h���\���" lP��R�*�BY4���x��{�;uK��4H|T��g)����Ά�з82K� H�R,?�q�X���F���s�!/e���u�w�̩ʷ��뷃�Y�S�5J��(�c�w�~S��ba��Ɗ3�