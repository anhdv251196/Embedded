XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��\~$t���Q�Mh�ģ	��>���)�T�:f��gU�*s��[7�q�:7��gn�ޅ MJߨ8aeԎ=�G�zb&�m��s�O�9��t�}�����̣���=���1�ƣ�Z��՘��;��j9�<Ֆ*���R3����ά�Ht��P�|E���`�'����N�3l��U.��>��fESZɵ�n'��HUy��v^|��@�u\X��$��Sz�B���c����1~� b�:��N�Ɉ�`^q�%4�t)�o��ӽOĂG2�W�9���b��$���7&D~e�u��/2��G�"�0Kc�5�'��9H!���q���"f���%^�����&OAD&ZS���%~�ۆF3he��s_�X�cxd��P����PiD�LX�=F\[[�O�OSa�u�v.('�n�.��Ō�%�Jfo���$�*�I�a{�ZeY^Лc.�~��sDٓ?��%�\p镙�0�OF��8�C��E��ˉ]�aZ8�`��C��C����ߐt����C�@M�n��^pO4���*�2;�$�Q�[��9p�j5�u�6���,�L:z&����2����l�*�����fd#j��l�-vQ��$}®7�_�1~QZ��x��?y����-Yk �l+��a���	
R��sy���g?����&n��&I�IPG�9�ъ�V��'��{�=a�Zk���1F��@.J<�ߗ���i��?��4�^���7��&��٫�ZI�ە�"��uLs��XlxVHYEB    1cf7     790Nѽ�?�oA���������;$+r�zi=��b[��}=�=����e'��u�?�y|���Ŭ�RV�i��C�_�;��F�#�5���w11^�AS�TJRL�\�͕����o> �����c�h��r-j3sOUv\��1�HZ���� �A�d6,�+�h���;ɥDn�mO��\��4( .#P(,:-��N�x �t_ܦ�+,3���nm���3�+H�Fh���[��#�<vX~��rk+Y��j�q5�闒�2[e�r�I��/� � "P��=�a'@��"��w֍3z�2����	RtD���c42����~H���*��<8^���u�^�A��.(��GSܩįv�,��g��v770?H��;�W8	aY�{�>��l�w�m���\$��PlC���8`���4����m˶A�!�)g�(uOe�e��ˉ��tI��!No�n�g�:�Tҋ#$���I	��QC`v}>J����A�n�ĳ$�KQ�zZ� ���Ap�p �p1�2$1Q�-k�٥ME��.1������`8k��ö���.+B���Sj��K�rf�c�iB>��{2�3
yz����ڔ�=\�b�(��&�O���O<�+5��9�
�&z���&ǂ�C�;�eJB��	��\P�q��ܑ�v�� D�����.�Y�0m��JC\걜Ž�-�ج���!��`�s���}���j]f�#K�dz��I�G�S�����d��X�z���=�����D�ҋ�rO��L߇���oJ���n����xu%N�������\�+��n����U&a�!��dGV>aj��hZ}�&���-������0���<!��Ks�CF�m��U�� fIDl�6)�Ix+�+�A?�D�c Z��=�q�`�C��rJ|�� 8N����UR��O2��38׮fo
�,�'���.5��[F<����hu�Ye�f�3��V�E�\ �]F�o�'"�^5e�T��,��9��G��D���w�a��0�>V	?��d�ʉH�!ǡA��g���գ�1�H��u�����{Ĺ�,ب8��W�u@�q��]+n��<H1^(
�[Ơ�s��4B�Ӕ64�"V�A��p�5Y����FJ��6��pi�o���6)�/5 p��H@�3<�	���z����K32@��}#J���G��Jo&���p�P_�%-<���6�_�����g'ݤjg{I^�[���)�cw��6���HQXd��wh
�M�@o�K���%\�MŠ)fiR�l3�Wkj��a��tb�&!��4��Z��w&���h�^x�-�8A=�'JKFZ�M�=�n��"ƙj}w6	��[��~�����'*��n}�QIn�f/L'��)-�ޢ2������Ǵ�F�{��ʛ5/��X��&�ǚ7���Ǉ�.��_d��2"K3 �΃ŷ�m��8��}l�A�6B[�ݾ3�����Ƅ�	�ޥ/`oQ�}���Z@-�t�\
�-R��>Ͼ�������x�S�� �'1ɸ�F��B�օ���>�{���׭#o�Vw^җ�i!���+}Rq�e�b�&�U@*�&՝�Șk��)�_`�k^���E�R��L�E�C>�-��8�9�`�R3lj���u�~k�]+֜��-��7�ц��p�J���v�
Ē벟�%�����
������y�}���w� �&g�Z����� [LOxbc�g��`Ss�����f:o��M;�lC@H�n;��W�$��b&Tr��3�5�",4x����߁���� ��*P�(����^�<�B)19W#�%a�хt_.>"u�^l�[ԟ��D�p�R�I�M�|��\������c_��#9
㫿pw�����W]�J�"u����K.W%O�L�æ�P�Tr����K����G�O�A�"