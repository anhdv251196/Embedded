XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��/k^kw�V�����K%@���-t�c��󼀚k��u9(QjR� ���Tn�B�d�� m܋ƄŪzܭ3��n-õ촰���4����c�jf��h0��!���<֕jSӢ5k�C�~&BkLii��83�+/����&i���Ș?�r��2v��Ɇ-��v��b�c���dDհ�����N4�_3�	�8ͬ �.c��RҺz ���G�s�z�@�3	]�Θ�.�<
2p��^J�Nh��׳7��ߟ���A�q<�`Vnv�6�|1�ɸbx0:v's_uz���-T��G ��=6��lRK!�$)��/�Ǌb��W &�W�8����Ά�=�M{K�9f������E��FA��9�Lg��Ž�f�	t���s�&m����xE�4�����i��<��ZR@W��s92���w����^�9-���^F�LxcGҒ%�^af8�қ٥�yɴQㆠk�C;U1'\�����Y�B��V���O���^a<n�A� ���
g\�-���=�f�g&�jJ�Ԁ2iQS����iZ�>+�#�!�A������ �*����L�Ϝ����Y/>���/��A��Cd���wȄ��MD9L�H%����N>�U���8[�il����W�S��+��Rw�/���f���7^X��_��E$DD4߹�(��wU�� �����F�E	'frRm�����}>���k�OG8k=n'�-�/.ؤ|wE�Q"�£s�%����Q!t�}���~�=��"���eE�{ �XlxVHYEB    1621     410��"�)�CbV�u�cƋ��q"ጤ]��a��@���$��1R�=mO�̀'���y8�.C�gc���`��
�b��[� 1�^*��3�u�n�I�A�&�h��'z�����4�~Z�czƗ���kHB�S��p'^��~���<��|9��c��V%Wad~�������J��z0��>r�>��0J��U��L�n��� �b�|��Z�[�Y�Sʦ��9�.c.����ӄ�a˷���S�\z�5���	�ӧ�,�NE��8x�O7�_�,�^Z�3k�����YEa��|��~Mx��`X��9~h�My�M��=�}�9=�Q���4p6�vB�ߥ���
�ёzT��$�N������<���Ȏ�R'���iyg��|!�ޤ���FZyʙ�V~��� �҈�Gr��(k޿Z��ҟz�pބ�f$%�CV��g�"��p�
�a0�>�ɯf����҄�l�/h�PR�;}�<��q?8�&�ۣ;�Cˋ�!�g%����N\�GJB�Tk���������I�Ǌ��(y��:Y~���\���bB���6�1�"�:7ۖ��Z���'�С����?ok�dGS�Ϣ^�0�L��6�:SQ<U���B�(���#����Wz0�T,�>.�2���y�sΗ�Ė;�	3��R�'D�$Tr���4����H�C�^[U��`e��{��),�M�v��DQG�������_(?�|��"����*�Q�<莩�Xٍ�AN��N�lW"����9�P� �͛%G^�Jm��@�N���Fq@2�Ƹ�}�IM��5"`d]�f���7���{�%Y>���	$5��8s5C��+�D��0���'Q��HX�y'��m�1�|S(�&E����>��U#�Z"�OM;W�P-ӨNE^(=#z5�:{;���F%	s�kj�`�k�	q�����l���o�TOAN�����i��q�\p��1gC8u�#$=���b����Rչ�:ZD��� #aU"XX�8�\�l�G��