XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���rV�Mg2G.���\�C -����wr2�e1���9��0Tw����n��St���y�*���"�4
�(�~u�QF�o�v,�b��A�ڑ�7�W�
�ʹ�/���)�0������/?f�^,w"����̝Y�Z�q�Nb��I�=h��Ifo�����������o�kG/��R�?o�s������onx�\�`7;���������D
aC�~�xΡ�Q���o#�\m�}�t�S�����~��s
�	���s���2x�ǔg*jV�y��"�n���L#)������&���g�S�m(Պ�;L$�qDr�Z�,����`�;��q*Dp.�i��7�S��\�#T��G7ʠ�4�hU
��8�ȴ��o��s
����+��M���7RfU&�R��:�����5_��ā��%)LM5,���������N�#>�H^�i���)�Z&�o�f�다CJ�}�qBi;��O�T�?Xi�����.0���`����kg�~BA���.�m���������K�(����Ŵ�,�^��$�-V��`�"��� CZ�S�u�3w)�lS�h��ޝ��0տ�tX�$[Y������D?:��0��M)�I�9`-��0A+S���j���-���5h�:�e	J�q}c���3>��&�e���.J�df�d��t
/u������H��?��"��� v(�#H[e�~Q���Aa�]��(�>��`1#+��W4&n� ��FOvXlxVHYEB    152d     580[qU���p��lT�̗_�g*&�
����*I���_o����|�+[�cu N�ֹ{90�U.��R����K�^C��&��)-ha��Y�M�����\��i!w�e�_��p{�YY4q�ID�ה�ypz���&�IVO���g2p��7�Ǻ8��yI�����rj�ҨxPlr�ؿ�X�(�	v�J�xœ'�L4�	#1��.7���i�Ee��j�ɵ@�Ӌn����]|��%��f�)�e��{���r��r��*���	�u��OF� *$��&�ۭ;C��0OPV���@,��)����o��"�
��=@��Tm�~��u0*���fk>^��b,+��j�F}]?V��O'�MT��b( U��џ�H�Z��g�X^�n9�$�u�r΄����P��E%66Y\���V�z�Rܠ�`H�jmu0�s���C]�f������UHNK����$:uև8įh�f��
�khQKY�6H�I���\0�w:0�&�����������(Փ�m�(MO��R��A�e��}]��=������]/��oI�K��e�= ȉ�~|�gB �wG���N��g�k��`/1�����J��09���0� �A����Em�}}�����/d�ش�[�/z��2 �3Ցe��"R�$R��.o��A�l�r��[ӕ�l-E������ͥ�3�L��J�/"��A���.!L�#)F���pzX��<D��	���f l���1u�R+��Ys��
���@����km�0��!���1y��6�� Lͅ� �e�*ɭ��O��$ZX%��d�@����R�r~�u!�X��ܯhF;��R��&������ ��-LװA�A��1��J��-�����
�ItI��mP7�I4�N�f�DD��B��K��qs���Oe#��5"Z�D�B���#FO|��ׄ��!��U�7j�U���x�P���CP�X^���R�eh�p^�7˙S��4L+��nm��ä��.y�ڿ�0�R��l�u<ވU�6���70��䡯�i�7M9��W�t�5�����)_�+��8�*w~>�����O{��s ����VN��4��̱�i�:���N�n��U��N{�2CrD����[��`�DY �4=�&��ņ&n\�{9-�+'���"J�BEG�6rm�B4�Y��S��ۊ� ����H�Yn���BQ�G��;���Gd:f�N�S�o�DVH�!�����b��J	k�A��I^ �6��;�u�3�y@�|��?~A-�x�?��6W���
���@#���֞բ��"���X��
^e;�+!� �+��Ћ�{�~��0�;����L*VNsZ>���,ሖ��<��n�������~����7Oֱ