XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���~��w/%]/PJ�J��ϭ��i�uL�-�3�7�r�Q����7�N��ƾ�K4����2-�z6=��0�|�Z�9R8P'.����>��Mj���_u�U8,���ͅ�9'�y����gP����D_��\�Hr��YO~�C5��8��7�n�� au.W@��f����g����3�>��^"?u���3��*$�&y4/�����t`�Г�)t��0�<j
Y��?���/�.�b�7�+{�� �{���R�?Q����g���1v��F�J����D1�����r���ΰ�;>PBUS	�3Zɾ��r��k+���}��x���S�J�(�Hu=����&�5����-T���$GN�;"�m+"��Ě��z�Ar���X�J3��V���4�t�����S�^nkK�j��D�x$WNS�LE�ր@B	�q�s��gg�sܱ�lJ[s��!�qƜ4| �T�@C�.��4�ݐ��)H�N��Rw�_?f A����-($✆������X��X>��'��Tr�_p*0>���x���������{9G��L'0�K�.����C����*!(��^��Kt��9(#���)<��;7�]�/\e����ƈbF#���Q��C= �8~�}������P�/��o�/����o���0�@5���=���I���d�x�� ɒ~�6ʔ*�<�9��@�@������,�M_T>;%kEl˄��B���B�SglY}p��SRm�L�����S�b����>^.A������XlxVHYEB    152b     580�[Q4��tni��@s��@uL\�s��zVe	Ģs䄎+h|�q�m����aB�$��	��'��(uy�P}54q8��^��sW���3�!��$�l6����XV+؂L��	kR�j����4�*��b{����Jhd�1�z;�̬�!����aq�aUl�8�5y(ˁ�uΣ����7�l��6-*��N�$i��2���qx���}��ӟ[�K�P�屌�YۗW
PmuOȜ��fUON�27���o��q�#K�����֬�5�fs�-�7��X�$y�i�H�����x7�[�p�
�RA���WKP�����U�ג�ǨV��&�	�w�SޑC�tǻ��S`���lk�GH�+b�1X�*�]rp3���Q{LƟ]�P����T.�H)B�1�vs1ԑI���'_x ,�4G�0V� �Ï��rm1�D�}L<t��K���(��A�N�����b>�ĥ�g�Z��\j����37�		`N-��X���(-��Xrq�p �nү���������.�i&»O�UL"�̺2Ŝ�v�����������M�0:�R��8+�<e=�R�дc��;��F|�c��8Y}��j��tz8`�p�h_>(ྒྷFs���H���"� %�.���A���o+?1�'�K!h��\�,���.Re��$��#fc�������t��������g�5Aڽ�X(�eGĝI���ȍ�a�W�_�,#_c�����kiZ����n�� (Pl`�ް��6�+2+UY�v���hPBr7��;Y+��Z�iC0�s���8@���>h�8�<��I�aќ�+��v������Y�-�u��N̗��u{��n�(������?׳ڻ�09Y\�gh�B�;��;� ��= ��������zY�l睕z65-P�L�K�Eg�7��\hj��1%}1MG�|��"�Kd{4h��_�f�9H���B{����gm����m�u�]����=��A%r��,���o\I����mQ���U�
*���&��#m��;G�a��e��5�2���9�{ɺ��D��יC�:z+���c�����K���V)ǰ�{
�:��BQkx��c#���b�-D�����W�>�~N�ǠW;�ߚ�X(�1t��c5�J��IS�,8�ڶ6S#ޮ�6�C�[�NQ�E�g�\%�}O������6���0��~���6{���T.%���A-B�
61z�8������4+=�.ˠr��4OO��"Rc�D����a�}9^���X�Z��FD	���n����� n0��H@2��R�"0^�k�/�P�g��O�s��~)gqn�KJr�S�ic#P��T_����o���8;2��r��^��9���%:9̟��4�ڐ� �D�<wc4�y�,��;��7"8�