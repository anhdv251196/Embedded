XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����.s�W���.�99��Ţ�q[Z3�����ݿDd�3���1P�]zn�qޮ�b+���I��	��*��K�\��@`��@ݯ�1����.&�L�S0��0,��8g���ќ?hH�,�|RhT�$�jP&u�ܗ�Dz���Ѕ{����}���Y�I,�?Х>$ȲG��z��gc_�ʶ:�呧 �i�
��K�a&�D�K�Np�����o+�P����
�8�s���w���U�%ݶ)LM�o����*�sCQ>vv�6g[1t1�w'��;��E��&�n�\Z�P�)�H�63�(ͰNuw+�<.y0�5�Da�3?�ߌ�]�&p;�lw8Q�Ӭk�4Np�ε*�lʹ�,ͱ��JK�'((������.]!�.�Bc}Ȁؔ��vt9��-�|<	d��:f��y��f<
�YCބ0"Gq��|/C��]���̚��1\�3Q�N���$	������� e�/���� c4���ְ;?�_�Rۗ*wv��棭ư-�LF���+Q����/5[g���c��fƣq蕳���u�Q߼Y�᫓�S�}��fjӹ�]�{��O�8��� `%����B� �H��4�F���tX�d�����C���~���L&��Ӑ[M3$)�^��9CQ��̕'?�a>�y�#)�d�Gv���=S���6$t@}�&(tq6��t����L�U����L ������:F�̀$H�߻U���Y
`��?u�0s���y	��9Z����)Ht���7|�`eE2B���u��7XlxVHYEB    41a2     c20��H�m6:V_�W��{�q$5O�Dd�WE�l���[8��p_C�/�j'� �/��-Q0԰=#W�āe�Հ�f8�I�Ͳ>��)���C���Tdnr��4e��q�]�4�ή-5�ڂ�A)�x-�&��c�����E�����Ǡ4�Իý����T�e��V�J`��ָPe���x��,1r,r?�Os��}Z�)�xp��߮���uؙy�g-]�L���d\1���̝�(\P�Fw����/�G��iZ�+��߸��0s�k�"��¢O�^� �H��B����s�[*ɪ�Ш,l�c�E\��Y�9y����,u�Z��^uD��f��J��7Z:r��I��]01H�
yn�����QD�w�!�}$�mR�s s�Cֆ]>��a��m6�1�-��DlLxf{wP�¦���,�՜�
M�fǣ8J�B�"����� �PCE�u�7a+C����㘨!ʾ��ߩ�z������N����Y�)�i��d�ʺ�c�;��a�5�ـ��[QkX0٥�u"���l�>{y4� jq��+_VA�j��S�u.�;�����7/��Z�zb�'���Q���f}p��C��{b1�]��3��3�/@�*޹�����6؜ �O���n+pj���I�I���>�c�xJ���13��/�Dc�{����(:�~�&��؄���|�wՈ�2�i9Mɲ��?��fjR��W��&/N~��! ��,��o���Iɳ�Х�}ju�ԅ�-Fn#�ϣB��O��$E��SWcCOM�}bc ���)��%o�%叻U��9��|٨��*C(B�j�s5��O���h���f%�����$�s�Ŷ!�b�ظ>��'ό�u���HtCM�"���f��kt �WNU�{�q�GB��{� �C" ���\�[�	�l�JU�����[����j0�j�+�C�mڹd�&�����9�K`x�@l�򩸦���j�����!Uva\�X)�����Z�=��]��`���D��T�/���F����� x�[�T)�9 6y�V�z�&6!��*LY͏��iE��-��:CQ��t�G歶0�N��w��s�\�Z��E����@�N�v1�-�+Q���'?��>/��t�l
�3T���/{Q�~6�r�ͳA����P��tb#���a
��M��'�F�박X�-�bl"�����ԕCQ�?�'�d�lx��
[z椿��ZgR��B�z����}�8d� c��JD���
zAK�j7J�a1u�����ZŪ���_�Z�L����uJո�n,q����� ������8+�	�����hS�s�����KM�a)kr���h���c��Koﴠ�$|@�eki�A�+��X+�=(*7{�EM,U��-�U�a����_�P�ܱ%�ڊyZ��wş9]�Sl��(�MKNG-d��jL�?�t=��#�9�\v=i2��bUǬ* �\�� ���Ky����TC�ə��o��s�7�>����0lHFE�a��� ww�z(9xV�n����`�RdP��@�5�(���m㤕�����>�W�����7�N��s̳�q5{wI�8����!%{ه��H�2�&sφͬv�kG?w��>������0���ǃx�	b2��Ԟ6ڡ�i#��@�y5Խ� �&x�]Qq���qic'P�^v�����걐�� y�f弲}jM����3)�
d��l}�˩�2��Jq�;�����i!���"��O����B:���$�>�]��Sa�`G% �(�u���_����;��0�ܝzǆ�u�?Kd�]�ݥ��I�-p�@�D�.��g�v�g�ۈ$�e8���e���{(�鶡��b�>2�N<�:�4�a,�B��q��-����3x5��3�FG1�j��Z'<!�����������tzu�;'����a���طH<��
�TH#��cN�@W���Gгv�R9�L{�	D&����S�N����w��@xH�2�3�{��yy��~�kv�������3�s��>�E؃=��!R@�d@٣",x�GL��t �� ��h�ȅ�Y�麈p��F�	�Q�	��7t��8P9���7m;���n1��cT%�F6�,vi߶�C�4!$��.��Jl����N����������-:���K	�<�Ȋ0�8}����SMd��K���GB���4�d�͑?����U���Oy'�|�	5�-�ܠ�>�gs!�1i���������WA�{���_�e �]u�ӛX��ʯ��R���4�%���&uI�����Z���m=v���� ݗ�k�;����S*�����\h�u��V{vQW��|�4#A���p��V
w�Ь��9����ᰬ��裺�\�o��4�ڞ��#a1&�W t ���Œ�;w���l���T�!ARC^���@ 9�N�/�c�ꕄΡ7M`\y뇗x'q�x�'x~��q�D��&t�l8Yvq��:��iD�y��^���N�:�۩���Tg���
;��jQ܌�u��}�����q��从z��dV��_�s��u��et���,r?� x�}�����/���8X���ɳ	HB�)���h�w@Ht�c��˟��$��^˾'����Xg���!�*���(�W�����Z�ؾ���5�i.3`���ڬˤ��zIZ�x��rL�M�3�1�5S���́%��V�Ϗ�˫l�y�:��<���xn9���;e�>Ԕ�;�o0�;��De���S��$�MhΪ��_ �����zލ�j%�.��X���v��ũl� ��.Cf�����d��$Ǒ�.�3� ��x$��1e)$�9R�A�x�AX���U9&������v�t|���Zs��Xjލ�yG��"6N�Ʒ�1s��c.��(r��S�i�y��cXpq[S5^��\?R�1�O��?���Ih�Y��Q������<�d��f.�k�lOc�� p�G$������B�J���8�{ռ���&q���<y�}�iLJ��f��\
�œJ�C։�<h"S�u�^��6�&(�*��>V