XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����Ȇ8w����U�+����4����Q�AC��E�����͸����ǺbA1�{�U8c\����GZ�IF#����d��f��0rpV�W E?k�=JX�������qA����x�'��;�!�dH��:K&���sE�����C������k�y���q9n^b'&�ˈa�r�!/�\�Z,?��H=�,Z̫�Gɔ4���e�E7��ABy1�Ҡ[�L����Mk�q�שz�b��.��b�9PZI1�d�@�$
�MQ)E����?�������~�6�S��(�0�'�� �ITP<�K�;�<=����:��,)���PčU�0��+&&Q�r@Y̤;�-�� �	�4W���8%h5A�A���~��U�<j�4v��F̀߁7�L����:��ⱙ*VD �e/ �|I��FDɫ�����.��8*��J��������e@�Zoܸ�x%`R��)U���5���ƽ���L���D��� �K����]�A��|@\\蕕t���U��V�v�qI*�ْr�O��$�_��QG�X>0���0��\H(Z���ٸ!�p>�.)ñ���wIs���V��݇=>���*�;��dN�<r�d�Ir�egR�0j�+��nة�ڌ]n�h����TBu��8��U\�FHa2�ؓ
�n��a�]�7���f�x�S!�4�-�QAg���C�imZ�uP]S�E1��vU�u�Qk�do
���O
�&�%�0�a�H�d�sr��OA��@������ϳ7	��ZXlxVHYEB    690c     b10�}���<70PDgw.�ĸ�k���@6��8��j�|���R.<TA�^N7�jf�Փ�����7�ix�7���e�g�xv1f�VU3���1�ף1"�����p9-矯���w��u�����r߂�ώv��f��ں���Lr�TM���>wu�w�}Мc8~�;5�/)N�iY��!y���� ����ͯ9q6�8]V��}���\ꞵ���Nܽ�5�&l���A�@�|�8�d� +R˒���a�*����n���m<։$c�`B�74��ɖ"9ԓ��+Յ��x�9����s��I��b�����^O-6�SC�%���l��1����/�6;���ӌ	�:D�����ގAY��ܣ_9��!C^\���ͺ-�����B�āth.�;xI�ui��6P ��aF1rg���k��f�BqK��aK����9��n�9�p1r�e�-w<L�,on�I�����GY@�)g����v\P|b�ƍ{�~[���w�z��U��� Ԗe�R!�N��!�3�:۾(D��NXB��'���$XLG�Ϸ�q�ȧ'X����[\�3Ff�0�>������N�Y�
Z����͒�Ӌ�b�����$�同>_ ���m�q��
>��3F�/�������0�3���Q2���#t�IH�^4\C	5�wG�:R���K�^���1��v|�xy0��i��˿�e�h0�y��Ռ�Q{��-����c��z�.��Lǅ2��GKu���G'�S��o���]b�S|?de7�vD"j��$��Ӳ�M]�)<�jv�g�^W�Vy;W���9�u��T4����W�Ș;t� i�/{ĕY�����\��(#���?�x��&�jK���J�z�6t�>�1�^���	����+"	�"����-q��-�<���;��ʔ��0���_�x��9� V��y���b:��"|QGj{5�F�yͦ�-b�r}�D�ߠ.�ش�����)�ي?
�6`���U��~`�=:# F�z���]0]�bJ�<�vxP���h�2��1�qu=�N��������x��Lm[��E����C����Zٮ���I����]%��==�,�E���Sr;NR��o(�貑6�����G͉���b��NȹC��#�,Gs�DH!�����w���:�i�pPMtA��fJ5�H�{�\U��N��'��3JroK>�u��x�U l=��8x"���� ��λ|�b�'2rNn��,ׂ[�/kr\�/�����
d�?D�k�-t�#�V����z ����n��&w��#AyK����ޘ�'�Ұ��E@Rdɞ�L�wXkW.71P�qB����S��&��m�fW��S��h��
$I�M�V��,{����������;�F��`i�<�%ț��Tv.^�,g�ϻ�ƽ���S@�����M�Ӊuȫ�%����z�S&�`Ѷ��B���@�Gr]Z݊V[�����싍<�C�F�Ϫ��y.��F�17t�ߖ�d�:#���@���`Z
W����J�a�-@�ԲWʇ���!A�iMd�o�#=���j����*J(��Q�V*��	"�r�30�T�{���ԆQ���ÛkET0���b����L��q��~T �S������l�cw�˭��2%�e�q��V�{!�*�;3um'Ne}=�c~��ع8�1O�w�xHH �8�aE��4�߸��I��k�a@҆�y,�K�C�b��Qp�/���� �<(���=z7˖��1���Iu��;��r}�a��k_��^.�ϭxV7�#e: �E���WcW��^`�YR�V\LsC�meez]��D"��3g%���Ő�l�nTȔ\Ph��:�n9�(-Q
�R ����\KK�`�C]�&*WC2y܉y��202u�r0�A�/�ĜP19pHG3�Y%{��3�Ơc&�	;�[�V]k��i��\�Ѐ29ߟ�>���K��ʣ2��"@~�ܹ�
���>��#�4����/vVtF\��#?���O�=�眞Bڱ8�����t1J�R�[������d���6�x�>g��D�{\0`�$7��N�e)�
=������T��y,~�c�ՕN�0��K���=�2w�zpZ��޲���,{ϵ����m�pϸ��4�A�U�`Ǟ1z4MYB����y;{[�s��a:\����m��u�d���'�Q:	��[1���p�tQ>�y�ŭ�:*V�p�W[LUIT)�U�$���2�SC�����S��|m	�t ��.k�x��r�5�w�p�xo��P_ED���q�m�F���A2c�$�i�Y:j2�(=���9�;2*���4���+L��YXLYFϭ\l��O�D���)�F���1�o�Zu�Љ��z�8|����]��JN��9eZ�kqE�=���ܥ5aDT֝��6�0�f�&2G�{"����&x��ǯ�7���n=��'M���%?�ܔ�t���X^p�Aau�E�C)li��=6+�`=2�:�����r	7L_��j����Ff�0:�����˾ڪ	��H�P+�b��J���d}����&�[4�WN�'Z�bl��Y��a�����2�cc����6�(H]6�]ƛD��x��60e���igl����"T�p�@Il�����j��+S��I�j(�LkUݧ�A��S���Y�n�`g����/U/p�k'_���R��i���(>�~�j��LS���d�=��7�n;���翐y���e|upF�f\����lE D���w����57�wˠ�����������2�3��*�H