XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��)���ض�N�-�b�S�v^�	:�U�r�����O���c4�g*a�5T�������v/v��Vr��M��Qc���=m��e��YE���I �Lk�..�������D�e)d�m
��N��H�����;�?e�C��������n�X۔��Y'�=�^��/�!�i�s�㾛�����I��63G���҄�1xJ�F.-�4�=):�3bpj|Z��A��,Н,Qd5Rr^���|$.s�?�Ӧ8blP�b�<����7ni�Ű噆�F\�J>h
ly01�_/.�ó�G �NQ*��O��֚��s�D�����ZX�j���P�$z�R�Q�(�*�vd1%���;ɊjP }��2_�����`�y��ih���2��'=D�&�-��*��H��Ϭ���CJO�ߓT]�����.!ϸD�wEu���|V]Q��kw�/V�f]��ݢ�m�6�\W��L�(n6$c:4��Ѫ�y��Li�d,Y�S=A;#Uȡ6��~
e:�]Ku���a�j�Gm2�,�'��8�#yX�J,�դPx�{��YicWm(����/�p��8����А��UB�������ت7F���āb}�}X�Ҡ�&����p	�2Π}�G�!��qh� s�g�"�S}Qyp�,8U��w}7�47T=���mγ���U7�i��\a����
��!?)^.Ά#MW$ܩ��j 'P�:xyS^��@p��Q�d�D�/!�/b�B��cw�ȦXlxVHYEB    1585     5b0�N}6�B8ڸ�q�]}+R�(�HSW��$�k��,G���r�y�Zf��+f�ф�5fdݬ���>�Q�����'Q���m��b���j	���.��́6(��p�hq�@6W[�����C���C�&��b���K1 �ỷfb-E{���gq|�������C�GL��+V!�x#u�/RP�^%�{J�,
d��?.��n�vfϻ�֒o��Y� �N��F뇎�_/�a�ƗC& Rɔ$[����"��㒀�/w�a9O0����f^}#�%�ЧUM�a�1��A��0v�fo8/ee]3n A� Q�~|�_��v*����H���ηm\oF�)�㓙z4�.I���Ԝ�K�n1-H^�anHVסg7��kd?��hW������������(����qqoR@����Z|�%�w��T�a�M�~*��+20�jA�R�8(U�.%c!���5�ze<4f�J߅A��5mKv7��t�蔣�{E��V3����||!�7X~pd9�%�ӌ��[|��P�Ss7h��ns|�C+e[O7�����霵=_��8־�L�n)5�m����ipNݽ�	���ƪ2��\UKLHΜ�oAbf&C~1�\�c����3���=+��p�����W��	�旡��||��IU����Aj�OG���D�TLzr�w�VYL��� ڢ��ڼ�l�[�!���}](�W��%a�D�hޮ9.
.E��w"2�-d	ף�-L�������7w'��w�Ne�?.�]�"ѓ>]^��/�X����Enq1����O�&a�{0cEOĈz��'F��!�9���2k9q�N�A~o�s��9�č���0W|�GF)L}�a"o� b&�{�{����Ax�k�ഀ�)\��yJ��I�[v'��x��O|d�Sm�
36%�R�������]q����Mp����MR��/��#�栺ГY(� ��)�)ws��GX�Np7�k�v8�òEm��� o�J,g�g��$�!GS�����ʌ�4,��\e��pA�~��cY�+�0��z2I����R*
f�����~'��4̬t;���dJ������]�aUC�"P6{��&�_��b�.tM�=��o��!M�:�?�|�n�uN1ά�B�c�^�W�0\�>t��G�!�%=�7Z�K��]%o����V�tA�� �ɥ,���L���h�����V,U�������K�{��+�j;���A��>#6}�r���HFS"JǊ+�I2Ӂ�i�-��Dp�*��[�e�Z�^aR����g��_�l�SJy|�w8�ՠ�6ɲ�+$���Kپ����,�N�B^��N=�"Vó�y���Xp1|@+�;�)i���)��D}z4[�"k�Qci��T�S�l��_��C��֌��q ���]ڲ�Y@a�İ�Xn
[�^x+`�|�l��0�=��b2�K��%